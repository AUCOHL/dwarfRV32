module rv32_CPU_v2 ( gnd!, vdd!, clk, rst, bdo, rfRS1, rfRS2, extR, extDone, IRQ, IRQnum, bdi, baddr, bsz, bwr, rfwr, rfrd, rfrs1, rfrs2, rfD, extA, extB, extStart, extFunc3);

input gnd!, vdd!;
input clk;
input rst;
input extDone;
input IRQ;
output bwr;
output rfwr;
output extStart;
input [31:0] bdo;
input [31:0] rfRS1;
input [31:0] rfRS2;
input [31:0] extR;
input [3:0] IRQnum;
output [31:0] bdi;
output [31:0] baddr;
output [1:0] bsz;
output [4:0] rfrd;
output [4:0] rfrs1;
output [4:0] rfrs2;
output [31:0] rfD;
output [31:0] extA;
output [31:0] extB;
output [2:0] extFunc3;

BUX2 BUX2_1 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_cyc_bF_buf8), .Q(CTRL_cyc_bF_buf0_bF_buf3) );
BUX2 BUX2_2 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_cyc_bF_buf14), .Q(CTRL_cyc_bF_buf0_bF_buf2) );
BUX2 BUX2_3 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_cyc_bF_buf4), .Q(CTRL_cyc_bF_buf0_bF_buf1) );
BUX2 BUX2_4 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_cyc_bF_buf0), .Q(CTRL_cyc_bF_buf0_bF_buf0) );
BUX2 BUX2_5 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_cyc_bF_buf8), .Q(CTRL_cyc_bF_buf1_bF_buf3) );
BUX2 BUX2_6 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_cyc_bF_buf1), .Q(CTRL_cyc_bF_buf1_bF_buf2) );
BUX2 BUX2_7 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_cyc_bF_buf13), .Q(CTRL_cyc_bF_buf1_bF_buf1) );
BUX2 BUX2_8 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_cyc_bF_buf2), .Q(CTRL_cyc_bF_buf1_bF_buf0) );
BUX2 BUX2_9 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_cyc_bF_buf2), .Q(CTRL_cyc_bF_buf2_bF_buf3) );
BUX2 BUX2_10 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_cyc_bF_buf3), .Q(CTRL_cyc_bF_buf2_bF_buf2) );
BUX2 BUX2_11 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_cyc_bF_buf7), .Q(CTRL_cyc_bF_buf2_bF_buf1) );
BUX2 BUX2_12 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_cyc_bF_buf2), .Q(CTRL_cyc_bF_buf2_bF_buf0) );
BUX2 BUX2_13 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_cyc_bF_buf3), .Q(CTRL_cyc_bF_buf3_bF_buf3) );
BUX2 BUX2_14 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_cyc_bF_buf11), .Q(CTRL_cyc_bF_buf3_bF_buf2) );
BUX2 BUX2_15 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_cyc_bF_buf13), .Q(CTRL_cyc_bF_buf3_bF_buf1) );
BUX2 BUX2_16 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_cyc_bF_buf0), .Q(CTRL_cyc_bF_buf3_bF_buf0) );
BUX2 BUX2_17 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_cyc_bF_buf9), .Q(CTRL_cyc_bF_buf4_bF_buf3) );
BUX2 BUX2_18 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_cyc_bF_buf4), .Q(CTRL_cyc_bF_buf4_bF_buf2) );
BUX2 BUX2_19 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_cyc_bF_buf5), .Q(CTRL_cyc_bF_buf4_bF_buf1) );
BUX2 BUX2_20 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_cyc_bF_buf4), .Q(CTRL_cyc_bF_buf4_bF_buf0) );
BUX2 BUX2_21 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_cyc_bF_buf0), .Q(CTRL_cyc_bF_buf5_bF_buf3) );
BUX2 BUX2_22 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_cyc_bF_buf10), .Q(CTRL_cyc_bF_buf5_bF_buf2) );
BUX2 BUX2_23 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_cyc_bF_buf4), .Q(CTRL_cyc_bF_buf5_bF_buf1) );
BUX2 BUX2_24 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_cyc_bF_buf5), .Q(CTRL_cyc_bF_buf5_bF_buf0) );
BUX2 BUX2_25 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_cyc_bF_buf6), .Q(CTRL_cyc_bF_buf6_bF_buf3) );
BUX2 BUX2_26 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_cyc_bF_buf3), .Q(CTRL_cyc_bF_buf6_bF_buf2) );
BUX2 BUX2_27 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_cyc_bF_buf7), .Q(CTRL_cyc_bF_buf6_bF_buf1) );
BUX2 BUX2_28 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_cyc_bF_buf6), .Q(CTRL_cyc_bF_buf6_bF_buf0) );
BUX2 BUX2_29 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_cyc_bF_buf7), .Q(CTRL_cyc_bF_buf7_bF_buf3) );
BUX2 BUX2_30 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_cyc_bF_buf12), .Q(CTRL_cyc_bF_buf7_bF_buf2) );
BUX2 BUX2_31 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_cyc_bF_buf7), .Q(CTRL_cyc_bF_buf7_bF_buf1) );
BUX2 BUX2_32 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_cyc_bF_buf5), .Q(CTRL_cyc_bF_buf7_bF_buf0) );
BUX2 BUX2_33 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_cyc_bF_buf8), .Q(CTRL_cyc_bF_buf8_bF_buf3) );
BUX2 BUX2_34 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_cyc_bF_buf1), .Q(CTRL_cyc_bF_buf8_bF_buf2) );
BUX2 BUX2_35 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_cyc_bF_buf5), .Q(CTRL_cyc_bF_buf8_bF_buf1) );
BUX2 BUX2_36 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_cyc_bF_buf11), .Q(CTRL_cyc_bF_buf8_bF_buf0) );
BUX2 BUX2_37 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_cyc_bF_buf4), .Q(CTRL_cyc_bF_buf9_bF_buf3) );
BUX2 BUX2_38 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_cyc_bF_buf9), .Q(CTRL_cyc_bF_buf9_bF_buf2) );
BUX2 BUX2_39 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_cyc_bF_buf2), .Q(CTRL_cyc_bF_buf9_bF_buf1) );
BUX2 BUX2_40 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_cyc_bF_buf14), .Q(CTRL_cyc_bF_buf9_bF_buf0) );
BUX2 BUX2_41 ( .gnd!(gnd!), .vdd!(vdd!), .A(clk), .Q(clk_hier0_bF_buf6) );
BUX2 BUX2_42 ( .gnd!(gnd!), .vdd!(vdd!), .A(clk), .Q(clk_hier0_bF_buf5) );
BUX2 BUX2_43 ( .gnd!(gnd!), .vdd!(vdd!), .A(clk), .Q(clk_hier0_bF_buf4) );
BUX2 BUX2_44 ( .gnd!(gnd!), .vdd!(vdd!), .A(clk), .Q(clk_hier0_bF_buf3) );
BUX2 BUX2_45 ( .gnd!(gnd!), .vdd!(vdd!), .A(clk), .Q(clk_hier0_bF_buf2) );
BUX2 BUX2_46 ( .gnd!(gnd!), .vdd!(vdd!), .A(clk), .Q(clk_hier0_bF_buf1) );
BUX2 BUX2_47 ( .gnd!(gnd!), .vdd!(vdd!), .A(clk), .Q(clk_hier0_bF_buf0) );
BUX2 BUX2_48 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_cyc_bF_buf1), .Q(CTRL_cyc_bF_buf10_bF_buf3) );
BUX2 BUX2_49 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_cyc_bF_buf14), .Q(CTRL_cyc_bF_buf10_bF_buf2) );
BUX2 BUX2_50 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_cyc_bF_buf10), .Q(CTRL_cyc_bF_buf10_bF_buf1) );
BUX2 BUX2_51 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_cyc_bF_buf10), .Q(CTRL_cyc_bF_buf10_bF_buf0) );
BUX2 BUX2_52 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_cyc_bF_buf11), .Q(CTRL_cyc_bF_buf11_bF_buf3) );
BUX2 BUX2_53 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_cyc_bF_buf3), .Q(CTRL_cyc_bF_buf11_bF_buf2) );
BUX2 BUX2_54 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_cyc_bF_buf12), .Q(CTRL_cyc_bF_buf11_bF_buf1) );
BUX2 BUX2_55 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_cyc_bF_buf1), .Q(CTRL_cyc_bF_buf11_bF_buf0) );
BUX2 BUX2_56 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_cyc_bF_buf6), .Q(CTRL_cyc_bF_buf12_bF_buf3) );
BUX2 BUX2_57 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_cyc_bF_buf11), .Q(CTRL_cyc_bF_buf12_bF_buf2) );
BUX2 BUX2_58 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_cyc_bF_buf2), .Q(CTRL_cyc_bF_buf12_bF_buf1) );
BUX2 BUX2_59 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_cyc_bF_buf7), .Q(CTRL_cyc_bF_buf12_bF_buf0) );
BUX2 BUX2_60 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_cyc_bF_buf6), .Q(CTRL_cyc_bF_buf13_bF_buf3) );
BUX2 BUX2_61 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_cyc_bF_buf9), .Q(CTRL_cyc_bF_buf13_bF_buf2) );
BUX2 BUX2_62 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_cyc_bF_buf10), .Q(CTRL_cyc_bF_buf13_bF_buf1) );
BUX2 BUX2_63 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_cyc_bF_buf13), .Q(CTRL_cyc_bF_buf13_bF_buf0) );
BUX2 BUX2_64 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_cyc_bF_buf13), .Q(CTRL_cyc_bF_buf14_bF_buf3) );
BUX2 BUX2_65 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_cyc_bF_buf12), .Q(CTRL_cyc_bF_buf14_bF_buf2) );
BUX2 BUX2_66 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_cyc_bF_buf0), .Q(CTRL_cyc_bF_buf14_bF_buf1) );
BUX2 BUX2_67 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_cyc_bF_buf10), .Q(CTRL_cyc_bF_buf14_bF_buf0) );
BUX2 BUX2_68 ( .gnd!(gnd!), .vdd!(vdd!), .A(_3247_), .Q(_3247__bF_buf4) );
BUX2 BUX2_69 ( .gnd!(gnd!), .vdd!(vdd!), .A(_3247_), .Q(_3247__bF_buf3) );
BUX2 BUX2_70 ( .gnd!(gnd!), .vdd!(vdd!), .A(_3247_), .Q(_3247__bF_buf2) );
BUX2 BUX2_71 ( .gnd!(gnd!), .vdd!(vdd!), .A(_3247_), .Q(_3247__bF_buf1) );
BUX2 BUX2_72 ( .gnd!(gnd!), .vdd!(vdd!), .A(_3247_), .Q(_3247__bF_buf0) );
BUX2 BUX2_73 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2650_), .Q(_2650__bF_buf7) );
BUX2 BUX2_74 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2650_), .Q(_2650__bF_buf6) );
BUX2 BUX2_75 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2650_), .Q(_2650__bF_buf5) );
BUX2 BUX2_76 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2650_), .Q(_2650__bF_buf4) );
BUX2 BUX2_77 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2650_), .Q(_2650__bF_buf3) );
BUX2 BUX2_78 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2650_), .Q(_2650__bF_buf2) );
BUX2 BUX2_79 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2650_), .Q(_2650__bF_buf1) );
BUX2 BUX2_80 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2650_), .Q(_2650__bF_buf0) );
BUX2 BUX2_81 ( .gnd!(gnd!), .vdd!(vdd!), .A(_3244_), .Q(_3244__bF_buf4) );
BUX2 BUX2_82 ( .gnd!(gnd!), .vdd!(vdd!), .A(_3244_), .Q(_3244__bF_buf3) );
BUX2 BUX2_83 ( .gnd!(gnd!), .vdd!(vdd!), .A(_3244_), .Q(_3244__bF_buf2) );
BUX2 BUX2_84 ( .gnd!(gnd!), .vdd!(vdd!), .A(_3244_), .Q(_3244__bF_buf1) );
BUX2 BUX2_85 ( .gnd!(gnd!), .vdd!(vdd!), .A(_3244_), .Q(_3244__bF_buf0) );
BUX2 BUX2_86 ( .gnd!(gnd!), .vdd!(vdd!), .A(EXT_type), .Q(EXT_type_bF_buf6) );
BUX2 BUX2_87 ( .gnd!(gnd!), .vdd!(vdd!), .A(EXT_type), .Q(EXT_type_bF_buf5) );
BUX2 BUX2_88 ( .gnd!(gnd!), .vdd!(vdd!), .A(EXT_type), .Q(EXT_type_bF_buf4) );
BUX2 BUX2_89 ( .gnd!(gnd!), .vdd!(vdd!), .A(EXT_type), .Q(EXT_type_bF_buf3) );
BUX2 BUX2_90 ( .gnd!(gnd!), .vdd!(vdd!), .A(EXT_type), .Q(EXT_type_bF_buf2) );
BUX2 BUX2_91 ( .gnd!(gnd!), .vdd!(vdd!), .A(EXT_type), .Q(EXT_type_bF_buf1) );
BUX2 BUX2_92 ( .gnd!(gnd!), .vdd!(vdd!), .A(EXT_type), .Q(EXT_type_bF_buf0) );
BUX2 BUX2_93 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2647_), .Q(_2647__bF_buf4) );
BUX2 BUX2_94 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2647_), .Q(_2647__bF_buf3) );
BUX2 BUX2_95 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2647_), .Q(_2647__bF_buf2) );
BUX2 BUX2_96 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2647_), .Q(_2647__bF_buf1) );
BUX2 BUX2_97 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2647_), .Q(_2647__bF_buf0) );
BUX2 BUX2_98 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_cu_ext_hold), .Q(CTRL_cu_ext_hold_bF_buf6) );
BUX2 BUX2_99 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_cu_ext_hold), .Q(CTRL_cu_ext_hold_bF_buf5) );
BUX2 BUX2_100 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_cu_ext_hold), .Q(CTRL_cu_ext_hold_bF_buf4) );
BUX2 BUX2_101 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_cu_ext_hold), .Q(CTRL_cu_ext_hold_bF_buf3) );
BUX2 BUX2_102 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_cu_ext_hold), .Q(CTRL_cu_ext_hold_bF_buf2) );
BUX2 BUX2_103 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_cu_ext_hold), .Q(CTRL_cu_ext_hold_bF_buf1) );
BUX2 BUX2_104 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_cu_ext_hold), .Q(CTRL_cu_ext_hold_bF_buf0) );
BUX2 BUX2_105 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_IDEC1_cu_custom_inst), .Q(CTRL_IDEC1_cu_custom_inst_bF_buf5) );
BUX2 BUX2_106 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_IDEC1_cu_custom_inst), .Q(CTRL_IDEC1_cu_custom_inst_bF_buf4) );
BUX2 BUX2_107 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_IDEC1_cu_custom_inst), .Q(CTRL_IDEC1_cu_custom_inst_bF_buf3) );
BUX2 BUX2_108 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_IDEC1_cu_custom_inst), .Q(CTRL_IDEC1_cu_custom_inst_bF_buf2) );
BUX2 BUX2_109 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_IDEC1_cu_custom_inst), .Q(CTRL_IDEC1_cu_custom_inst_bF_buf1) );
BUX2 BUX2_110 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_IDEC1_cu_custom_inst), .Q(CTRL_IDEC1_cu_custom_inst_bF_buf0) );
BUX2 BUX2_111 ( .gnd!(gnd!), .vdd!(vdd!), .A(_682__0_), .Q(_682__0_bF_buf3) );
BUX2 BUX2_112 ( .gnd!(gnd!), .vdd!(vdd!), .A(_682__0_), .Q(_682__0_bF_buf2) );
BUX2 BUX2_113 ( .gnd!(gnd!), .vdd!(vdd!), .A(_682__0_), .Q(_682__0_bF_buf1) );
BUX2 BUX2_114 ( .gnd!(gnd!), .vdd!(vdd!), .A(_682__0_), .Q(_682__0_bF_buf0) );
BUX2 BUX2_115 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1242_), .Q(_1242__bF_buf4) );
BUX2 BUX2_116 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1242_), .Q(_1242__bF_buf3) );
BUX2 BUX2_117 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1242_), .Q(_1242__bF_buf2) );
BUX2 BUX2_118 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1242_), .Q(_1242__bF_buf1) );
BUX2 BUX2_119 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1242_), .Q(_1242__bF_buf0) );
BUX2 BUX2_120 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_cu_r2_src), .Q(CTRL_cu_r2_src_bF_buf5) );
BUX2 BUX2_121 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_cu_r2_src), .Q(CTRL_cu_r2_src_bF_buf4) );
BUX2 BUX2_122 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_cu_r2_src), .Q(CTRL_cu_r2_src_bF_buf3) );
BUX2 BUX2_123 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_cu_r2_src), .Q(CTRL_cu_r2_src_bF_buf2) );
BUX2 BUX2_124 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_cu_r2_src), .Q(CTRL_cu_r2_src_bF_buf1) );
BUX2 BUX2_125 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_cu_r2_src), .Q(CTRL_cu_r2_src_bF_buf0) );
BUX2 BUX2_126 ( .gnd!(gnd!), .vdd!(vdd!), .A(_476_), .Q(_476__bF_buf4) );
BUX2 BUX2_127 ( .gnd!(gnd!), .vdd!(vdd!), .A(_476_), .Q(_476__bF_buf3) );
BUX2 BUX2_128 ( .gnd!(gnd!), .vdd!(vdd!), .A(_476_), .Q(_476__bF_buf2) );
BUX2 BUX2_129 ( .gnd!(gnd!), .vdd!(vdd!), .A(_476_), .Q(_476__bF_buf1) );
BUX2 BUX2_130 ( .gnd!(gnd!), .vdd!(vdd!), .A(_476_), .Q(_476__bF_buf0) );
BUX2 BUX2_131 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1048_), .Q(_1048__bF_buf4) );
BUX2 BUX2_132 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1048_), .Q(_1048__bF_buf3) );
BUX2 BUX2_133 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1048_), .Q(_1048__bF_buf2) );
BUX2 BUX2_134 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1048_), .Q(_1048__bF_buf1) );
BUX2 BUX2_135 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1048_), .Q(_1048__bF_buf0) );
BUX2 BUX2_136 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_IDEC1_cu_load_inst), .Q(CTRL_IDEC1_cu_load_inst_bF_buf4) );
BUX2 BUX2_137 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_IDEC1_cu_load_inst), .Q(CTRL_IDEC1_cu_load_inst_bF_buf3) );
BUX2 BUX2_138 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_IDEC1_cu_load_inst), .Q(CTRL_IDEC1_cu_load_inst_bF_buf2) );
BUX2 BUX2_139 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_IDEC1_cu_load_inst), .Q(CTRL_IDEC1_cu_load_inst_bF_buf1) );
BUX2 BUX2_140 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_IDEC1_cu_load_inst), .Q(CTRL_IDEC1_cu_load_inst_bF_buf0) );
BUX2 BUX2_141 ( .gnd!(gnd!), .vdd!(vdd!), .A(_39_), .Q(_39__bF_buf4) );
BUX2 BUX2_142 ( .gnd!(gnd!), .vdd!(vdd!), .A(_39_), .Q(_39__bF_buf3) );
BUX2 BUX2_143 ( .gnd!(gnd!), .vdd!(vdd!), .A(_39_), .Q(_39__bF_buf2) );
BUX2 BUX2_144 ( .gnd!(gnd!), .vdd!(vdd!), .A(_39_), .Q(_39__bF_buf1) );
BUX2 BUX2_145 ( .gnd!(gnd!), .vdd!(vdd!), .A(_39_), .Q(_39__bF_buf0) );
BUX2 BUX2_146 ( .gnd!(gnd!), .vdd!(vdd!), .A(_952_), .Q(_952__bF_buf5) );
BUX2 BUX2_147 ( .gnd!(gnd!), .vdd!(vdd!), .A(_952_), .Q(_952__bF_buf4) );
BUX2 BUX2_148 ( .gnd!(gnd!), .vdd!(vdd!), .A(_952_), .Q(_952__bF_buf3) );
BUX2 BUX2_149 ( .gnd!(gnd!), .vdd!(vdd!), .A(_952_), .Q(_952__bF_buf2) );
BUX2 BUX2_150 ( .gnd!(gnd!), .vdd!(vdd!), .A(_952_), .Q(_952__bF_buf1) );
BUX2 BUX2_151 ( .gnd!(gnd!), .vdd!(vdd!), .A(_952_), .Q(_952__bF_buf0) );
BUX2 BUX2_152 ( .gnd!(gnd!), .vdd!(vdd!), .A(clk_hier0_bF_buf5), .Q(clk_bF_buf53) );
BUX2 BUX2_153 ( .gnd!(gnd!), .vdd!(vdd!), .A(clk_hier0_bF_buf0), .Q(clk_bF_buf52) );
BUX2 BUX2_154 ( .gnd!(gnd!), .vdd!(vdd!), .A(clk_hier0_bF_buf2), .Q(clk_bF_buf51) );
BUX2 BUX2_155 ( .gnd!(gnd!), .vdd!(vdd!), .A(clk_hier0_bF_buf3), .Q(clk_bF_buf50) );
BUX2 BUX2_156 ( .gnd!(gnd!), .vdd!(vdd!), .A(clk_hier0_bF_buf2), .Q(clk_bF_buf49) );
BUX2 BUX2_157 ( .gnd!(gnd!), .vdd!(vdd!), .A(clk_hier0_bF_buf0), .Q(clk_bF_buf48) );
BUX2 BUX2_158 ( .gnd!(gnd!), .vdd!(vdd!), .A(clk_hier0_bF_buf6), .Q(clk_bF_buf47) );
BUX2 BUX2_159 ( .gnd!(gnd!), .vdd!(vdd!), .A(clk_hier0_bF_buf4), .Q(clk_bF_buf46) );
BUX2 BUX2_160 ( .gnd!(gnd!), .vdd!(vdd!), .A(clk_hier0_bF_buf1), .Q(clk_bF_buf45) );
BUX2 BUX2_161 ( .gnd!(gnd!), .vdd!(vdd!), .A(clk_hier0_bF_buf1), .Q(clk_bF_buf44) );
BUX2 BUX2_162 ( .gnd!(gnd!), .vdd!(vdd!), .A(clk_hier0_bF_buf1), .Q(clk_bF_buf43) );
BUX2 BUX2_163 ( .gnd!(gnd!), .vdd!(vdd!), .A(clk_hier0_bF_buf3), .Q(clk_bF_buf42) );
BUX2 BUX2_164 ( .gnd!(gnd!), .vdd!(vdd!), .A(clk_hier0_bF_buf3), .Q(clk_bF_buf41) );
BUX2 BUX2_165 ( .gnd!(gnd!), .vdd!(vdd!), .A(clk_hier0_bF_buf4), .Q(clk_bF_buf40) );
BUX2 BUX2_166 ( .gnd!(gnd!), .vdd!(vdd!), .A(clk_hier0_bF_buf1), .Q(clk_bF_buf39) );
BUX2 BUX2_167 ( .gnd!(gnd!), .vdd!(vdd!), .A(clk_hier0_bF_buf2), .Q(clk_bF_buf38) );
BUX2 BUX2_168 ( .gnd!(gnd!), .vdd!(vdd!), .A(clk_hier0_bF_buf6), .Q(clk_bF_buf37) );
BUX2 BUX2_169 ( .gnd!(gnd!), .vdd!(vdd!), .A(clk_hier0_bF_buf5), .Q(clk_bF_buf36) );
BUX2 BUX2_170 ( .gnd!(gnd!), .vdd!(vdd!), .A(clk_hier0_bF_buf0), .Q(clk_bF_buf35) );
BUX2 BUX2_171 ( .gnd!(gnd!), .vdd!(vdd!), .A(clk_hier0_bF_buf3), .Q(clk_bF_buf34) );
BUX2 BUX2_172 ( .gnd!(gnd!), .vdd!(vdd!), .A(clk_hier0_bF_buf1), .Q(clk_bF_buf33) );
BUX2 BUX2_173 ( .gnd!(gnd!), .vdd!(vdd!), .A(clk_hier0_bF_buf4), .Q(clk_bF_buf32) );
BUX2 BUX2_174 ( .gnd!(gnd!), .vdd!(vdd!), .A(clk_hier0_bF_buf3), .Q(clk_bF_buf31) );
BUX2 BUX2_175 ( .gnd!(gnd!), .vdd!(vdd!), .A(clk_hier0_bF_buf3), .Q(clk_bF_buf30) );
BUX2 BUX2_176 ( .gnd!(gnd!), .vdd!(vdd!), .A(clk_hier0_bF_buf3), .Q(clk_bF_buf29) );
BUX2 BUX2_177 ( .gnd!(gnd!), .vdd!(vdd!), .A(clk_hier0_bF_buf4), .Q(clk_bF_buf28) );
BUX2 BUX2_178 ( .gnd!(gnd!), .vdd!(vdd!), .A(clk_hier0_bF_buf6), .Q(clk_bF_buf27) );
BUX2 BUX2_179 ( .gnd!(gnd!), .vdd!(vdd!), .A(clk_hier0_bF_buf4), .Q(clk_bF_buf26) );
BUX2 BUX2_180 ( .gnd!(gnd!), .vdd!(vdd!), .A(clk_hier0_bF_buf2), .Q(clk_bF_buf25) );
BUX2 BUX2_181 ( .gnd!(gnd!), .vdd!(vdd!), .A(clk_hier0_bF_buf1), .Q(clk_bF_buf24) );
BUX2 BUX2_182 ( .gnd!(gnd!), .vdd!(vdd!), .A(clk_hier0_bF_buf4), .Q(clk_bF_buf23) );
BUX2 BUX2_183 ( .gnd!(gnd!), .vdd!(vdd!), .A(clk_hier0_bF_buf5), .Q(clk_bF_buf22) );
BUX2 BUX2_184 ( .gnd!(gnd!), .vdd!(vdd!), .A(clk_hier0_bF_buf5), .Q(clk_bF_buf21) );
BUX2 BUX2_185 ( .gnd!(gnd!), .vdd!(vdd!), .A(clk_hier0_bF_buf0), .Q(clk_bF_buf20) );
BUX2 BUX2_186 ( .gnd!(gnd!), .vdd!(vdd!), .A(clk_hier0_bF_buf5), .Q(clk_bF_buf19) );
BUX2 BUX2_187 ( .gnd!(gnd!), .vdd!(vdd!), .A(clk_hier0_bF_buf0), .Q(clk_bF_buf18) );
BUX2 BUX2_188 ( .gnd!(gnd!), .vdd!(vdd!), .A(clk_hier0_bF_buf6), .Q(clk_bF_buf17) );
BUX2 BUX2_189 ( .gnd!(gnd!), .vdd!(vdd!), .A(clk_hier0_bF_buf0), .Q(clk_bF_buf16) );
BUX2 BUX2_190 ( .gnd!(gnd!), .vdd!(vdd!), .A(clk_hier0_bF_buf2), .Q(clk_bF_buf15) );
BUX2 BUX2_191 ( .gnd!(gnd!), .vdd!(vdd!), .A(clk_hier0_bF_buf5), .Q(clk_bF_buf14) );
BUX2 BUX2_192 ( .gnd!(gnd!), .vdd!(vdd!), .A(clk_hier0_bF_buf6), .Q(clk_bF_buf13) );
BUX2 BUX2_193 ( .gnd!(gnd!), .vdd!(vdd!), .A(clk_hier0_bF_buf4), .Q(clk_bF_buf12) );
BUX2 BUX2_194 ( .gnd!(gnd!), .vdd!(vdd!), .A(clk_hier0_bF_buf6), .Q(clk_bF_buf11) );
BUX2 BUX2_195 ( .gnd!(gnd!), .vdd!(vdd!), .A(clk_hier0_bF_buf5), .Q(clk_bF_buf10) );
BUX2 BUX2_196 ( .gnd!(gnd!), .vdd!(vdd!), .A(clk_hier0_bF_buf1), .Q(clk_bF_buf9) );
BUX2 BUX2_197 ( .gnd!(gnd!), .vdd!(vdd!), .A(clk_hier0_bF_buf2), .Q(clk_bF_buf8) );
BUX2 BUX2_198 ( .gnd!(gnd!), .vdd!(vdd!), .A(clk_hier0_bF_buf5), .Q(clk_bF_buf7) );
BUX2 BUX2_199 ( .gnd!(gnd!), .vdd!(vdd!), .A(clk_hier0_bF_buf6), .Q(clk_bF_buf6) );
BUX2 BUX2_200 ( .gnd!(gnd!), .vdd!(vdd!), .A(clk_hier0_bF_buf6), .Q(clk_bF_buf5) );
BUX2 BUX2_201 ( .gnd!(gnd!), .vdd!(vdd!), .A(clk_hier0_bF_buf2), .Q(clk_bF_buf4) );
BUX2 BUX2_202 ( .gnd!(gnd!), .vdd!(vdd!), .A(clk_hier0_bF_buf2), .Q(clk_bF_buf3) );
BUX2 BUX2_203 ( .gnd!(gnd!), .vdd!(vdd!), .A(clk_hier0_bF_buf3), .Q(clk_bF_buf2) );
BUX2 BUX2_204 ( .gnd!(gnd!), .vdd!(vdd!), .A(clk_hier0_bF_buf4), .Q(clk_bF_buf1) );
BUX2 BUX2_205 ( .gnd!(gnd!), .vdd!(vdd!), .A(clk_hier0_bF_buf0), .Q(clk_bF_buf0) );
BUX2 BUX2_206 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1524_), .Q(_1524__bF_buf3) );
BUX2 BUX2_207 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1524_), .Q(_1524__bF_buf2) );
BUX2 BUX2_208 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1524_), .Q(_1524__bF_buf1) );
BUX2 BUX2_209 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1524_), .Q(_1524__bF_buf0) );
BUX2 BUX2_210 ( .gnd!(gnd!), .vdd!(vdd!), .A(_473_), .Q(_473__bF_buf5) );
BUX2 BUX2_211 ( .gnd!(gnd!), .vdd!(vdd!), .A(_473_), .Q(_473__bF_buf4) );
BUX2 BUX2_212 ( .gnd!(gnd!), .vdd!(vdd!), .A(_473_), .Q(_473__bF_buf3) );
BUX2 BUX2_213 ( .gnd!(gnd!), .vdd!(vdd!), .A(_473_), .Q(_473__bF_buf2) );
BUX2 BUX2_214 ( .gnd!(gnd!), .vdd!(vdd!), .A(_473_), .Q(_473__bF_buf1) );
BUX2 BUX2_215 ( .gnd!(gnd!), .vdd!(vdd!), .A(_473_), .Q(_473__bF_buf0) );
BUX2 BUX2_216 ( .gnd!(gnd!), .vdd!(vdd!), .A(CNTR_ld_cycle), .Q(CNTR_ld_cycle_bF_buf6) );
BUX2 BUX2_217 ( .gnd!(gnd!), .vdd!(vdd!), .A(CNTR_ld_cycle), .Q(CNTR_ld_cycle_bF_buf5) );
BUX2 BUX2_218 ( .gnd!(gnd!), .vdd!(vdd!), .A(CNTR_ld_cycle), .Q(CNTR_ld_cycle_bF_buf4) );
BUX2 BUX2_219 ( .gnd!(gnd!), .vdd!(vdd!), .A(CNTR_ld_cycle), .Q(CNTR_ld_cycle_bF_buf3) );
BUX2 BUX2_220 ( .gnd!(gnd!), .vdd!(vdd!), .A(CNTR_ld_cycle), .Q(CNTR_ld_cycle_bF_buf2) );
BUX2 BUX2_221 ( .gnd!(gnd!), .vdd!(vdd!), .A(CNTR_ld_cycle), .Q(CNTR_ld_cycle_bF_buf1) );
BUX2 BUX2_222 ( .gnd!(gnd!), .vdd!(vdd!), .A(CNTR_ld_cycle), .Q(CNTR_ld_cycle_bF_buf0) );
BUX2 BUX2_223 ( .gnd!(gnd!), .vdd!(vdd!), .A(_36_), .Q(_36__bF_buf3) );
BUX2 BUX2_224 ( .gnd!(gnd!), .vdd!(vdd!), .A(_36_), .Q(_36__bF_buf2) );
BUX2 BUX2_225 ( .gnd!(gnd!), .vdd!(vdd!), .A(_36_), .Q(_36__bF_buf1) );
BUX2 BUX2_226 ( .gnd!(gnd!), .vdd!(vdd!), .A(_36_), .Q(_36__bF_buf0) );
BUX2 BUX2_227 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1233_), .Q(_1233__bF_buf4) );
BUX2 BUX2_228 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1233_), .Q(_1233__bF_buf3) );
BUX2 BUX2_229 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1233_), .Q(_1233__bF_buf2) );
BUX2 BUX2_230 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1233_), .Q(_1233__bF_buf1) );
BUX2 BUX2_231 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1233_), .Q(_1233__bF_buf0) );
BUX2 BUX2_232 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1230_), .Q(_1230__bF_buf5) );
BUX2 BUX2_233 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1230_), .Q(_1230__bF_buf4) );
BUX2 BUX2_234 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1230_), .Q(_1230__bF_buf3) );
BUX2 BUX2_235 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1230_), .Q(_1230__bF_buf2) );
BUX2 BUX2_236 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1230_), .Q(_1230__bF_buf1) );
BUX2 BUX2_237 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1230_), .Q(_1230__bF_buf0) );
BUX2 BUX2_238 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1227_), .Q(_1227__bF_buf6) );
BUX2 BUX2_239 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1227_), .Q(_1227__bF_buf5) );
BUX2 BUX2_240 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1227_), .Q(_1227__bF_buf4) );
BUX2 BUX2_241 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1227_), .Q(_1227__bF_buf3) );
BUX2 BUX2_242 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1227_), .Q(_1227__bF_buf2) );
BUX2 BUX2_243 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1227_), .Q(_1227__bF_buf1) );
BUX2 BUX2_244 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1227_), .Q(_1227__bF_buf0) );
BUX2 BUX2_245 ( .gnd!(gnd!), .vdd!(vdd!), .A(_3117_), .Q(_3117__bF_buf7) );
BUX2 BUX2_246 ( .gnd!(gnd!), .vdd!(vdd!), .A(_3117_), .Q(_3117__bF_buf6) );
BUX2 BUX2_247 ( .gnd!(gnd!), .vdd!(vdd!), .A(_3117_), .Q(_3117__bF_buf5) );
BUX2 BUX2_248 ( .gnd!(gnd!), .vdd!(vdd!), .A(_3117_), .Q(_3117__bF_buf4) );
BUX2 BUX2_249 ( .gnd!(gnd!), .vdd!(vdd!), .A(_3117_), .Q(_3117__bF_buf3) );
BUX2 BUX2_250 ( .gnd!(gnd!), .vdd!(vdd!), .A(_3117_), .Q(_3117__bF_buf2) );
BUX2 BUX2_251 ( .gnd!(gnd!), .vdd!(vdd!), .A(_3117_), .Q(_3117__bF_buf1) );
BUX2 BUX2_252 ( .gnd!(gnd!), .vdd!(vdd!), .A(_3117_), .Q(_3117__bF_buf0) );
BUX2 BUX2_253 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1221_), .Q(_1221__bF_buf4) );
BUX2 BUX2_254 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1221_), .Q(_1221__bF_buf3) );
BUX2 BUX2_255 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1221_), .Q(_1221__bF_buf2) );
BUX2 BUX2_256 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1221_), .Q(_1221__bF_buf1) );
BUX2 BUX2_257 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1221_), .Q(_1221__bF_buf0) );
BUX2 BUX2_258 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2329_), .Q(_2329__bF_buf4) );
BUX2 BUX2_259 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2329_), .Q(_2329__bF_buf3) );
BUX2 BUX2_260 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2329_), .Q(_2329__bF_buf2) );
BUX2 BUX2_261 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2329_), .Q(_2329__bF_buf1) );
BUX2 BUX2_262 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2329_), .Q(_2329__bF_buf0) );
BUX2 BUX2_263 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2367_), .Q(_2367__bF_buf4) );
BUX2 BUX2_264 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2367_), .Q(_2367__bF_buf3) );
BUX2 BUX2_265 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2367_), .Q(_2367__bF_buf2) );
BUX2 BUX2_266 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2367_), .Q(_2367__bF_buf1) );
BUX2 BUX2_267 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2367_), .Q(_2367__bF_buf0) );
BUX2 BUX2_268 ( .gnd!(gnd!), .vdd!(vdd!), .A(_21_), .Q(_21__bF_buf7) );
BUX2 BUX2_269 ( .gnd!(gnd!), .vdd!(vdd!), .A(_21_), .Q(_21__bF_buf6) );
BUX2 BUX2_270 ( .gnd!(gnd!), .vdd!(vdd!), .A(_21_), .Q(_21__bF_buf5) );
BUX2 BUX2_271 ( .gnd!(gnd!), .vdd!(vdd!), .A(_21_), .Q(_21__bF_buf4) );
BUX2 BUX2_272 ( .gnd!(gnd!), .vdd!(vdd!), .A(_21_), .Q(_21__bF_buf3) );
BUX2 BUX2_273 ( .gnd!(gnd!), .vdd!(vdd!), .A(_21_), .Q(_21__bF_buf2) );
BUX2 BUX2_274 ( .gnd!(gnd!), .vdd!(vdd!), .A(_21_), .Q(_21__bF_buf1) );
BUX2 BUX2_275 ( .gnd!(gnd!), .vdd!(vdd!), .A(_21_), .Q(_21__bF_buf0) );
BUX2 BUX2_276 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_cu_r1_src), .Q(CTRL_cu_r1_src_bF_buf3) );
BUX2 BUX2_277 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_cu_r1_src), .Q(CTRL_cu_r1_src_bF_buf2) );
BUX2 BUX2_278 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_cu_r1_src), .Q(CTRL_cu_r1_src_bF_buf1) );
BUX2 BUX2_279 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_cu_r1_src), .Q(CTRL_cu_r1_src_bF_buf0) );
BUX2 BUX2_280 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_IDEC1_cu_system_inst), .Q(CTRL_IDEC1_cu_system_inst_bF_buf7) );
BUX2 BUX2_281 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_IDEC1_cu_system_inst), .Q(CTRL_IDEC1_cu_system_inst_bF_buf6) );
BUX2 BUX2_282 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_IDEC1_cu_system_inst), .Q(CTRL_IDEC1_cu_system_inst_bF_buf5) );
BUX2 BUX2_283 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_IDEC1_cu_system_inst), .Q(CTRL_IDEC1_cu_system_inst_bF_buf4) );
BUX2 BUX2_284 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_IDEC1_cu_system_inst), .Q(CTRL_IDEC1_cu_system_inst_bF_buf3) );
BUX2 BUX2_285 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_IDEC1_cu_system_inst), .Q(CTRL_IDEC1_cu_system_inst_bF_buf2) );
BUX2 BUX2_286 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_IDEC1_cu_system_inst), .Q(CTRL_IDEC1_cu_system_inst_bF_buf1) );
BUX2 BUX2_287 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_IDEC1_cu_system_inst), .Q(CTRL_IDEC1_cu_system_inst_bF_buf0) );
BUX2 BUX2_288 ( .gnd!(gnd!), .vdd!(vdd!), .A(_931_), .Q(_931__bF_buf5) );
BUX2 BUX2_289 ( .gnd!(gnd!), .vdd!(vdd!), .A(_931_), .Q(_931__bF_buf4) );
BUX2 BUX2_290 ( .gnd!(gnd!), .vdd!(vdd!), .A(_931_), .Q(_931__bF_buf3) );
BUX2 BUX2_291 ( .gnd!(gnd!), .vdd!(vdd!), .A(_931_), .Q(_931__bF_buf2) );
BUX2 BUX2_292 ( .gnd!(gnd!), .vdd!(vdd!), .A(_931_), .Q(_931__bF_buf1) );
BUX2 BUX2_293 ( .gnd!(gnd!), .vdd!(vdd!), .A(_931_), .Q(_931__bF_buf0) );
BUX2 BUX2_294 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_cu_alu_b_src), .Q(CTRL_cu_alu_b_src_bF_buf4) );
BUX2 BUX2_295 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_cu_alu_b_src), .Q(CTRL_cu_alu_b_src_bF_buf3) );
BUX2 BUX2_296 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_cu_alu_b_src), .Q(CTRL_cu_alu_b_src_bF_buf2) );
BUX2 BUX2_297 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_cu_alu_b_src), .Q(CTRL_cu_alu_b_src_bF_buf1) );
BUX2 BUX2_298 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_cu_alu_b_src), .Q(CTRL_cu_alu_b_src_bF_buf0) );
BUX2 BUX2_299 ( .gnd!(gnd!), .vdd!(vdd!), .A(_3246_), .Q(_3246__bF_buf4) );
BUX2 BUX2_300 ( .gnd!(gnd!), .vdd!(vdd!), .A(_3246_), .Q(_3246__bF_buf3) );
BUX2 BUX2_301 ( .gnd!(gnd!), .vdd!(vdd!), .A(_3246_), .Q(_3246__bF_buf2) );
BUX2 BUX2_302 ( .gnd!(gnd!), .vdd!(vdd!), .A(_3246_), .Q(_3246__bF_buf1) );
BUX2 BUX2_303 ( .gnd!(gnd!), .vdd!(vdd!), .A(_3246_), .Q(_3246__bF_buf0) );
BUX2 BUX2_304 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2458_), .Q(_2458__bF_buf5) );
BUX2 BUX2_305 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2458_), .Q(_2458__bF_buf4) );
BUX2 BUX2_306 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2458_), .Q(_2458__bF_buf3) );
BUX2 BUX2_307 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2458_), .Q(_2458__bF_buf2) );
BUX2 BUX2_308 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2458_), .Q(_2458__bF_buf1) );
BUX2 BUX2_309 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2458_), .Q(_2458__bF_buf0) );
BUX2 BUX2_310 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1059_), .Q(_1059__bF_buf3) );
BUX2 BUX2_311 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1059_), .Q(_1059__bF_buf2) );
BUX2 BUX2_312 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1059_), .Q(_1059__bF_buf1) );
BUX2 BUX2_313 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1059_), .Q(_1059__bF_buf0) );
BUX2 BUX2_314 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1212_), .Q(_1212__bF_buf4) );
BUX2 BUX2_315 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1212_), .Q(_1212__bF_buf3) );
BUX2 BUX2_316 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1212_), .Q(_1212__bF_buf2) );
BUX2 BUX2_317 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1212_), .Q(_1212__bF_buf1) );
BUX2 BUX2_318 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1212_), .Q(_1212__bF_buf0) );
BUX2 BUX2_319 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2646_), .Q(_2646__bF_buf3) );
BUX2 BUX2_320 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2646_), .Q(_2646__bF_buf2) );
BUX2 BUX2_321 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2646_), .Q(_2646__bF_buf1) );
BUX2 BUX2_322 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2646_), .Q(_2646__bF_buf0) );
BUX2 BUX2_323 ( .gnd!(gnd!), .vdd!(vdd!), .A(_866_), .Q(_866__bF_buf5) );
BUX2 BUX2_324 ( .gnd!(gnd!), .vdd!(vdd!), .A(_866_), .Q(_866__bF_buf4) );
BUX2 BUX2_325 ( .gnd!(gnd!), .vdd!(vdd!), .A(_866_), .Q(_866__bF_buf3) );
BUX2 BUX2_326 ( .gnd!(gnd!), .vdd!(vdd!), .A(_866_), .Q(_866__bF_buf2) );
BUX2 BUX2_327 ( .gnd!(gnd!), .vdd!(vdd!), .A(_866_), .Q(_866__bF_buf1) );
BUX2 BUX2_328 ( .gnd!(gnd!), .vdd!(vdd!), .A(_866_), .Q(_866__bF_buf0) );
BUX2 BUX2_329 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2643_), .Q(_2643__bF_buf5) );
BUX2 BUX2_330 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2643_), .Q(_2643__bF_buf4) );
BUX2 BUX2_331 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2643_), .Q(_2643__bF_buf3) );
BUX2 BUX2_332 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2643_), .Q(_2643__bF_buf2) );
BUX2 BUX2_333 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2643_), .Q(_2643__bF_buf1) );
BUX2 BUX2_334 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2643_), .Q(_2643__bF_buf0) );
BUX2 BUX2_335 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_IDEC1_cu_auipc_inst), .Q(CTRL_IDEC1_cu_auipc_inst_bF_buf4) );
BUX2 BUX2_336 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_IDEC1_cu_auipc_inst), .Q(CTRL_IDEC1_cu_auipc_inst_bF_buf3) );
BUX2 BUX2_337 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_IDEC1_cu_auipc_inst), .Q(CTRL_IDEC1_cu_auipc_inst_bF_buf2) );
BUX2 BUX2_338 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_IDEC1_cu_auipc_inst), .Q(CTRL_IDEC1_cu_auipc_inst_bF_buf1) );
BUX2 BUX2_339 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_IDEC1_cu_auipc_inst), .Q(CTRL_IDEC1_cu_auipc_inst_bF_buf0) );
BUX2 BUX2_340 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_cu_csr_rd_s1), .Q(CTRL_cu_csr_rd_s1_bF_buf7) );
BUX2 BUX2_341 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_cu_csr_rd_s1), .Q(CTRL_cu_csr_rd_s1_bF_buf6) );
BUX2 BUX2_342 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_cu_csr_rd_s1), .Q(CTRL_cu_csr_rd_s1_bF_buf5) );
BUX2 BUX2_343 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_cu_csr_rd_s1), .Q(CTRL_cu_csr_rd_s1_bF_buf4) );
BUX2 BUX2_344 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_cu_csr_rd_s1), .Q(CTRL_cu_csr_rd_s1_bF_buf3) );
BUX2 BUX2_345 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_cu_csr_rd_s1), .Q(CTRL_cu_csr_rd_s1_bF_buf2) );
BUX2 BUX2_346 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_cu_csr_rd_s1), .Q(CTRL_cu_csr_rd_s1_bF_buf1) );
BUX2 BUX2_347 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_cu_csr_rd_s1), .Q(CTRL_cu_csr_rd_s1_bF_buf0) );
BUX2 BUX2_348 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1203_), .Q(_1203__bF_buf4) );
BUX2 BUX2_349 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1203_), .Q(_1203__bF_buf3) );
BUX2 BUX2_350 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1203_), .Q(_1203__bF_buf2) );
BUX2 BUX2_351 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1203_), .Q(_1203__bF_buf1) );
BUX2 BUX2_352 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1203_), .Q(_1203__bF_buf0) );
BUX2 BUX2_353 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1526_), .Q(_1526__bF_buf4) );
BUX2 BUX2_354 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1526_), .Q(_1526__bF_buf3) );
BUX2 BUX2_355 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1526_), .Q(_1526__bF_buf2) );
BUX2 BUX2_356 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1526_), .Q(_1526__bF_buf1) );
BUX2 BUX2_357 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1526_), .Q(_1526__bF_buf0) );
BUX2 BUX2_358 ( .gnd!(gnd!), .vdd!(vdd!), .A(_434_), .Q(_434__bF_buf3) );
BUX2 BUX2_359 ( .gnd!(gnd!), .vdd!(vdd!), .A(_434_), .Q(_434__bF_buf2) );
BUX2 BUX2_360 ( .gnd!(gnd!), .vdd!(vdd!), .A(_434_), .Q(_434__bF_buf1) );
BUX2 BUX2_361 ( .gnd!(gnd!), .vdd!(vdd!), .A(_434_), .Q(_434__bF_buf0) );
BUX2 BUX2_362 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1235_), .Q(_1235__bF_buf4) );
BUX2 BUX2_363 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1235_), .Q(_1235__bF_buf3) );
BUX2 BUX2_364 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1235_), .Q(_1235__bF_buf2) );
BUX2 BUX2_365 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1235_), .Q(_1235__bF_buf1) );
BUX2 BUX2_366 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1235_), .Q(_1235__bF_buf0) );
BUX2 BUX2_367 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1329_), .Q(_1329__bF_buf4) );
BUX2 BUX2_368 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1329_), .Q(_1329__bF_buf3) );
BUX2 BUX2_369 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1329_), .Q(_1329__bF_buf2) );
BUX2 BUX2_370 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1329_), .Q(_1329__bF_buf1) );
BUX2 BUX2_371 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1329_), .Q(_1329__bF_buf0) );
BUX2 BUX2_372 ( .gnd!(gnd!), .vdd!(vdd!), .A(_32_), .Q(_32__bF_buf4) );
BUX2 BUX2_373 ( .gnd!(gnd!), .vdd!(vdd!), .A(_32_), .Q(_32__bF_buf3) );
BUX2 BUX2_374 ( .gnd!(gnd!), .vdd!(vdd!), .A(_32_), .Q(_32__bF_buf2) );
BUX2 BUX2_375 ( .gnd!(gnd!), .vdd!(vdd!), .A(_32_), .Q(_32__bF_buf1) );
BUX2 BUX2_376 ( .gnd!(gnd!), .vdd!(vdd!), .A(_32_), .Q(_32__bF_buf0) );
BUX2 BUX2_377 ( .gnd!(gnd!), .vdd!(vdd!), .A(_29_), .Q(_29__bF_buf6) );
BUX2 BUX2_378 ( .gnd!(gnd!), .vdd!(vdd!), .A(_29_), .Q(_29__bF_buf5) );
BUX2 BUX2_379 ( .gnd!(gnd!), .vdd!(vdd!), .A(_29_), .Q(_29__bF_buf4) );
BUX2 BUX2_380 ( .gnd!(gnd!), .vdd!(vdd!), .A(_29_), .Q(_29__bF_buf3) );
BUX2 BUX2_381 ( .gnd!(gnd!), .vdd!(vdd!), .A(_29_), .Q(_29__bF_buf2) );
BUX2 BUX2_382 ( .gnd!(gnd!), .vdd!(vdd!), .A(_29_), .Q(_29__bF_buf1) );
BUX2 BUX2_383 ( .gnd!(gnd!), .vdd!(vdd!), .A(_29_), .Q(_29__bF_buf0) );
BUX2 BUX2_384 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2243_), .Q(_2243__bF_buf7) );
BUX2 BUX2_385 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2243_), .Q(_2243__bF_buf6) );
BUX2 BUX2_386 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2243_), .Q(_2243__bF_buf5) );
BUX2 BUX2_387 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2243_), .Q(_2243__bF_buf4) );
BUX2 BUX2_388 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2243_), .Q(_2243__bF_buf3) );
BUX2 BUX2_389 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2243_), .Q(_2243__bF_buf2) );
BUX2 BUX2_390 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2243_), .Q(_2243__bF_buf1) );
BUX2 BUX2_391 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2243_), .Q(_2243__bF_buf0) );
BUX2 BUX2_392 ( .gnd!(gnd!), .vdd!(vdd!), .A(CNTR_ld_timer), .Q(CNTR_ld_timer_bF_buf4) );
BUX2 BUX2_393 ( .gnd!(gnd!), .vdd!(vdd!), .A(CNTR_ld_timer), .Q(CNTR_ld_timer_bF_buf3) );
BUX2 BUX2_394 ( .gnd!(gnd!), .vdd!(vdd!), .A(CNTR_ld_timer), .Q(CNTR_ld_timer_bF_buf2) );
BUX2 BUX2_395 ( .gnd!(gnd!), .vdd!(vdd!), .A(CNTR_ld_timer), .Q(CNTR_ld_timer_bF_buf1) );
BUX2 BUX2_396 ( .gnd!(gnd!), .vdd!(vdd!), .A(CNTR_ld_timer), .Q(CNTR_ld_timer_bF_buf0) );
BUX2 BUX2_397 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1226_), .Q(_1226__bF_buf6) );
BUX2 BUX2_398 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1226_), .Q(_1226__bF_buf5) );
BUX2 BUX2_399 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1226_), .Q(_1226__bF_buf4) );
BUX2 BUX2_400 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1226_), .Q(_1226__bF_buf3) );
BUX2 BUX2_401 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1226_), .Q(_1226__bF_buf2) );
BUX2 BUX2_402 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1226_), .Q(_1226__bF_buf1) );
BUX2 BUX2_403 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1226_), .Q(_1226__bF_buf0) );
BUX2 BUX2_404 ( .gnd!(gnd!), .vdd!(vdd!), .A(_595_), .Q(_595__bF_buf4) );
BUX2 BUX2_405 ( .gnd!(gnd!), .vdd!(vdd!), .A(_595_), .Q(_595__bF_buf3) );
BUX2 BUX2_406 ( .gnd!(gnd!), .vdd!(vdd!), .A(_595_), .Q(_595__bF_buf2) );
BUX2 BUX2_407 ( .gnd!(gnd!), .vdd!(vdd!), .A(_595_), .Q(_595__bF_buf1) );
BUX2 BUX2_408 ( .gnd!(gnd!), .vdd!(vdd!), .A(_595_), .Q(_595__bF_buf0) );
BUX2 BUX2_409 ( .gnd!(gnd!), .vdd!(vdd!), .A(_23_), .Q(_23__bF_buf6) );
BUX2 BUX2_410 ( .gnd!(gnd!), .vdd!(vdd!), .A(_23_), .Q(_23__bF_buf5) );
BUX2 BUX2_411 ( .gnd!(gnd!), .vdd!(vdd!), .A(_23_), .Q(_23__bF_buf4) );
BUX2 BUX2_412 ( .gnd!(gnd!), .vdd!(vdd!), .A(_23_), .Q(_23__bF_buf3) );
BUX2 BUX2_413 ( .gnd!(gnd!), .vdd!(vdd!), .A(_23_), .Q(_23__bF_buf2) );
BUX2 BUX2_414 ( .gnd!(gnd!), .vdd!(vdd!), .A(_23_), .Q(_23__bF_buf1) );
BUX2 BUX2_415 ( .gnd!(gnd!), .vdd!(vdd!), .A(_23_), .Q(_23__bF_buf0) );
BUX2 BUX2_416 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_IDEC1_cu_jalr_inst), .Q(CTRL_IDEC1_cu_jalr_inst_bF_buf5) );
BUX2 BUX2_417 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_IDEC1_cu_jalr_inst), .Q(CTRL_IDEC1_cu_jalr_inst_bF_buf4) );
BUX2 BUX2_418 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_IDEC1_cu_jalr_inst), .Q(CTRL_IDEC1_cu_jalr_inst_bF_buf3) );
BUX2 BUX2_419 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_IDEC1_cu_jalr_inst), .Q(CTRL_IDEC1_cu_jalr_inst_bF_buf2) );
BUX2 BUX2_420 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_IDEC1_cu_jalr_inst), .Q(CTRL_IDEC1_cu_jalr_inst_bF_buf1) );
BUX2 BUX2_421 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_IDEC1_cu_jalr_inst), .Q(CTRL_IDEC1_cu_jalr_inst_bF_buf0) );
BUX2 BUX2_422 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1252_), .Q(_1252__bF_buf5) );
BUX2 BUX2_423 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1252_), .Q(_1252__bF_buf4) );
BUX2 BUX2_424 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1252_), .Q(_1252__bF_buf3) );
BUX2 BUX2_425 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1252_), .Q(_1252__bF_buf2) );
BUX2 BUX2_426 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1252_), .Q(_1252__bF_buf1) );
BUX2 BUX2_427 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1252_), .Q(_1252__bF_buf0) );
BUX2 BUX2_428 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2686_), .Q(_2686__bF_buf3) );
BUX2 BUX2_429 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2686_), .Q(_2686__bF_buf2) );
BUX2 BUX2_430 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2686_), .Q(_2686__bF_buf1) );
BUX2 BUX2_431 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2686_), .Q(_2686__bF_buf0) );
BUX2 BUX2_432 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_cu_pc_s2), .Q(CTRL_cu_pc_s2_bF_buf7) );
BUX2 BUX2_433 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_cu_pc_s2), .Q(CTRL_cu_pc_s2_bF_buf6) );
BUX2 BUX2_434 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_cu_pc_s2), .Q(CTRL_cu_pc_s2_bF_buf5) );
BUX2 BUX2_435 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_cu_pc_s2), .Q(CTRL_cu_pc_s2_bF_buf4) );
BUX2 BUX2_436 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_cu_pc_s2), .Q(CTRL_cu_pc_s2_bF_buf3) );
BUX2 BUX2_437 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_cu_pc_s2), .Q(CTRL_cu_pc_s2_bF_buf2) );
BUX2 BUX2_438 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_cu_pc_s2), .Q(CTRL_cu_pc_s2_bF_buf1) );
BUX2 BUX2_439 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_cu_pc_s2), .Q(CTRL_cu_pc_s2_bF_buf0) );
BUX2 BUX2_440 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_cu_pc_s3), .Q(CTRL_cu_pc_s3_bF_buf4) );
BUX2 BUX2_441 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_cu_pc_s3), .Q(CTRL_cu_pc_s3_bF_buf3) );
BUX2 BUX2_442 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_cu_pc_s3), .Q(CTRL_cu_pc_s3_bF_buf2) );
BUX2 BUX2_443 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_cu_pc_s3), .Q(CTRL_cu_pc_s3_bF_buf1) );
BUX2 BUX2_444 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_cu_pc_s3), .Q(CTRL_cu_pc_s3_bF_buf0) );
BUX2 BUX2_445 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_cu_pc_s4), .Q(CTRL_cu_pc_s4_bF_buf5) );
BUX2 BUX2_446 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_cu_pc_s4), .Q(CTRL_cu_pc_s4_bF_buf4) );
BUX2 BUX2_447 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_cu_pc_s4), .Q(CTRL_cu_pc_s4_bF_buf3) );
BUX2 BUX2_448 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_cu_pc_s4), .Q(CTRL_cu_pc_s4_bF_buf2) );
BUX2 BUX2_449 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_cu_pc_s4), .Q(CTRL_cu_pc_s4_bF_buf1) );
BUX2 BUX2_450 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_cu_pc_s4), .Q(CTRL_cu_pc_s4_bF_buf0) );
BUX2 BUX2_451 ( .gnd!(gnd!), .vdd!(vdd!), .A(_682__1_), .Q(_682__1_bF_buf4) );
BUX2 BUX2_452 ( .gnd!(gnd!), .vdd!(vdd!), .A(_682__1_), .Q(_682__1_bF_buf3) );
BUX2 BUX2_453 ( .gnd!(gnd!), .vdd!(vdd!), .A(_682__1_), .Q(_682__1_bF_buf2) );
BUX2 BUX2_454 ( .gnd!(gnd!), .vdd!(vdd!), .A(_682__1_), .Q(_682__1_bF_buf1) );
BUX2 BUX2_455 ( .gnd!(gnd!), .vdd!(vdd!), .A(_682__1_), .Q(_682__1_bF_buf0) );
BUX2 BUX2_456 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1240_), .Q(_1240__bF_buf6) );
BUX2 BUX2_457 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1240_), .Q(_1240__bF_buf5) );
BUX2 BUX2_458 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1240_), .Q(_1240__bF_buf4) );
BUX2 BUX2_459 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1240_), .Q(_1240__bF_buf3) );
BUX2 BUX2_460 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1240_), .Q(_1240__bF_buf2) );
BUX2 BUX2_461 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1240_), .Q(_1240__bF_buf1) );
BUX2 BUX2_462 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1240_), .Q(_1240__bF_buf0) );
BUX2 BUX2_463 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_cyc), .Q(CTRL_cyc_bF_buf14) );
BUX2 BUX2_464 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_cyc), .Q(CTRL_cyc_bF_buf13) );
BUX2 BUX2_465 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_cyc), .Q(CTRL_cyc_bF_buf12) );
BUX2 BUX2_466 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_cyc), .Q(CTRL_cyc_bF_buf11) );
BUX2 BUX2_467 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_cyc), .Q(CTRL_cyc_bF_buf10) );
BUX2 BUX2_468 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_cyc), .Q(CTRL_cyc_bF_buf9) );
BUX2 BUX2_469 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_cyc), .Q(CTRL_cyc_bF_buf8) );
BUX2 BUX2_470 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_cyc), .Q(CTRL_cyc_bF_buf7) );
BUX2 BUX2_471 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_cyc), .Q(CTRL_cyc_bF_buf6) );
BUX2 BUX2_472 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_cyc), .Q(CTRL_cyc_bF_buf5) );
BUX2 BUX2_473 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_cyc), .Q(CTRL_cyc_bF_buf4) );
BUX2 BUX2_474 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_cyc), .Q(CTRL_cyc_bF_buf3) );
BUX2 BUX2_475 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_cyc), .Q(CTRL_cyc_bF_buf2) );
BUX2 BUX2_476 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_cyc), .Q(CTRL_cyc_bF_buf1) );
BUX2 BUX2_477 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_cyc), .Q(CTRL_cyc_bF_buf0) );
BUX2 BUX2_478 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1525_), .Q(_1525__bF_buf4) );
BUX2 BUX2_479 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1525_), .Q(_1525__bF_buf3) );
BUX2 BUX2_480 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1525_), .Q(_1525__bF_buf2) );
BUX2 BUX2_481 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1525_), .Q(_1525__bF_buf1) );
BUX2 BUX2_482 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1525_), .Q(_1525__bF_buf0) );
BUX2 BUX2_483 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1143_), .Q(_1143__bF_buf4) );
BUX2 BUX2_484 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1143_), .Q(_1143__bF_buf3) );
BUX2 BUX2_485 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1143_), .Q(_1143__bF_buf2) );
BUX2 BUX2_486 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1143_), .Q(_1143__bF_buf1) );
BUX2 BUX2_487 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1143_), .Q(_1143__bF_buf0) );
BUX2 BUX2_488 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2195_), .Q(_2195__bF_buf3) );
BUX2 BUX2_489 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2195_), .Q(_2195__bF_buf2) );
BUX2 BUX2_490 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2195_), .Q(_2195__bF_buf1) );
BUX2 BUX2_491 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2195_), .Q(_2195__bF_buf0) );
BUX2 BUX2_492 ( .gnd!(gnd!), .vdd!(vdd!), .A(_909_), .Q(_909__bF_buf4) );
BUX2 BUX2_493 ( .gnd!(gnd!), .vdd!(vdd!), .A(_909_), .Q(_909__bF_buf3) );
BUX2 BUX2_494 ( .gnd!(gnd!), .vdd!(vdd!), .A(_909_), .Q(_909__bF_buf2) );
BUX2 BUX2_495 ( .gnd!(gnd!), .vdd!(vdd!), .A(_909_), .Q(_909__bF_buf1) );
BUX2 BUX2_496 ( .gnd!(gnd!), .vdd!(vdd!), .A(_909_), .Q(_909__bF_buf0) );
BUX2 BUX2_497 ( .gnd!(gnd!), .vdd!(vdd!), .A(_471_), .Q(_471__bF_buf7) );
BUX2 BUX2_498 ( .gnd!(gnd!), .vdd!(vdd!), .A(_471_), .Q(_471__bF_buf6) );
BUX2 BUX2_499 ( .gnd!(gnd!), .vdd!(vdd!), .A(_471_), .Q(_471__bF_buf5) );
BUX2 BUX2_500 ( .gnd!(gnd!), .vdd!(vdd!), .A(_471_), .Q(_471__bF_buf4) );
BUX2 BUX2_501 ( .gnd!(gnd!), .vdd!(vdd!), .A(_471_), .Q(_471__bF_buf3) );
BUX2 BUX2_502 ( .gnd!(gnd!), .vdd!(vdd!), .A(_471_), .Q(_471__bF_buf2) );
BUX2 BUX2_503 ( .gnd!(gnd!), .vdd!(vdd!), .A(_471_), .Q(_471__bF_buf1) );
BUX2 BUX2_504 ( .gnd!(gnd!), .vdd!(vdd!), .A(_471_), .Q(_471__bF_buf0) );
BUX2 BUX2_505 ( .gnd!(gnd!), .vdd!(vdd!), .A(ALU_func7_5_), .Q(ALU_func7_5_bF_buf3) );
BUX2 BUX2_506 ( .gnd!(gnd!), .vdd!(vdd!), .A(ALU_func7_5_), .Q(ALU_func7_5_bF_buf2) );
BUX2 BUX2_507 ( .gnd!(gnd!), .vdd!(vdd!), .A(ALU_func7_5_), .Q(ALU_func7_5_bF_buf1) );
BUX2 BUX2_508 ( .gnd!(gnd!), .vdd!(vdd!), .A(ALU_func7_5_), .Q(ALU_func7_5_bF_buf0) );
BUX2 BUX2_509 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1328_), .Q(_1328__bF_buf4) );
BUX2 BUX2_510 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1328_), .Q(_1328__bF_buf3) );
BUX2 BUX2_511 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1328_), .Q(_1328__bF_buf2) );
BUX2 BUX2_512 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1328_), .Q(_1328__bF_buf1) );
BUX2 BUX2_513 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1328_), .Q(_1328__bF_buf0) );
BUX2 BUX2_514 ( .gnd!(gnd!), .vdd!(vdd!), .A(_888_), .Q(_888__bF_buf4) );
BUX2 BUX2_515 ( .gnd!(gnd!), .vdd!(vdd!), .A(_888_), .Q(_888__bF_buf3) );
BUX2 BUX2_516 ( .gnd!(gnd!), .vdd!(vdd!), .A(_888_), .Q(_888__bF_buf2) );
BUX2 BUX2_517 ( .gnd!(gnd!), .vdd!(vdd!), .A(_888_), .Q(_888__bF_buf1) );
BUX2 BUX2_518 ( .gnd!(gnd!), .vdd!(vdd!), .A(_888_), .Q(_888__bF_buf0) );
BUX2 BUX2_519 ( .gnd!(gnd!), .vdd!(vdd!), .A(_941_), .Q(_941__bF_buf4) );
BUX2 BUX2_520 ( .gnd!(gnd!), .vdd!(vdd!), .A(_941_), .Q(_941__bF_buf3) );
BUX2 BUX2_521 ( .gnd!(gnd!), .vdd!(vdd!), .A(_941_), .Q(_941__bF_buf2) );
BUX2 BUX2_522 ( .gnd!(gnd!), .vdd!(vdd!), .A(_941_), .Q(_941__bF_buf1) );
BUX2 BUX2_523 ( .gnd!(gnd!), .vdd!(vdd!), .A(_941_), .Q(_941__bF_buf0) );
BUX2 BUX2_524 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1322_), .Q(_1322__bF_buf3) );
BUX2 BUX2_525 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1322_), .Q(_1322__bF_buf2) );
BUX2 BUX2_526 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1322_), .Q(_1322__bF_buf1) );
BUX2 BUX2_527 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1322_), .Q(_1322__bF_buf0) );
BUX2 BUX2_528 ( .gnd!(gnd!), .vdd!(vdd!), .A(_268_), .Q(_268__bF_buf8) );
BUX2 BUX2_529 ( .gnd!(gnd!), .vdd!(vdd!), .A(_268_), .Q(_268__bF_buf7) );
BUX2 BUX2_530 ( .gnd!(gnd!), .vdd!(vdd!), .A(_268_), .Q(_268__bF_buf6) );
BUX2 BUX2_531 ( .gnd!(gnd!), .vdd!(vdd!), .A(_268_), .Q(_268__bF_buf5) );
BUX2 BUX2_532 ( .gnd!(gnd!), .vdd!(vdd!), .A(_268_), .Q(_268__bF_buf4) );
BUX2 BUX2_533 ( .gnd!(gnd!), .vdd!(vdd!), .A(_268_), .Q(_268__bF_buf3) );
BUX2 BUX2_534 ( .gnd!(gnd!), .vdd!(vdd!), .A(_268_), .Q(_268__bF_buf2) );
BUX2 BUX2_535 ( .gnd!(gnd!), .vdd!(vdd!), .A(_268_), .Q(_268__bF_buf1) );
BUX2 BUX2_536 ( .gnd!(gnd!), .vdd!(vdd!), .A(_268_), .Q(_268__bF_buf0) );
BUX2 BUX2_537 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2371_), .Q(_2371__bF_buf3) );
BUX2 BUX2_538 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2371_), .Q(_2371__bF_buf2) );
BUX2 BUX2_539 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2371_), .Q(_2371__bF_buf1) );
BUX2 BUX2_540 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2371_), .Q(_2371__bF_buf0) );
BUX2 BUX2_541 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1222_), .Q(_1222__bF_buf5) );
BUX2 BUX2_542 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1222_), .Q(_1222__bF_buf4) );
BUX2 BUX2_543 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1222_), .Q(_1222__bF_buf3) );
BUX2 BUX2_544 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1222_), .Q(_1222__bF_buf2) );
BUX2 BUX2_545 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1222_), .Q(_1222__bF_buf1) );
BUX2 BUX2_546 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1222_), .Q(_1222__bF_buf0) );
NA2X1 NA2X1_1 ( .gnd!(gnd!), .vdd!(vdd!), .A(R_0_), .B(CTRL_cyc_bF_buf14_bF_buf0), .Q(_593_) );
NO2X1 NO2X1_1 ( .gnd!(gnd!), .vdd!(vdd!), .A(ALU_r_0_), .B(CTRL_IDEC1_cu_custom_inst_bF_buf5), .Q(_594_) );
INX2 INX2_1 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_IDEC1_cu_custom_inst_bF_buf3), .Q(_595_) );
NO2X1 NO2X1_2 ( .gnd!(gnd!), .vdd!(vdd!), .A(extR[0]), .B(_595__bF_buf2), .Q(_596_) );
ON31X1 ON31X1_1 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_cyc_bF_buf13_bF_buf1), .B(_594_), .C(_596_), .D(_593_), .Q(_6__0_) );
NA2X1 NA2X1_2 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_cyc_bF_buf12_bF_buf0), .B(R_1_), .Q(_597_) );
NO2X1 NO2X1_3 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_IDEC1_cu_custom_inst_bF_buf0), .B(ALU_r_1_), .Q(_598_) );
NO2X1 NO2X1_4 ( .gnd!(gnd!), .vdd!(vdd!), .A(extR[1]), .B(_595__bF_buf2), .Q(_599_) );
ON31X1 ON31X1_2 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_cyc_bF_buf11_bF_buf3), .B(_598_), .C(_599_), .D(_597_), .Q(_6__1_) );
NA2X1 NA2X1_3 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_cyc_bF_buf10_bF_buf3), .B(R_2_), .Q(_600_) );
NO2X1 NO2X1_5 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_IDEC1_cu_custom_inst_bF_buf2), .B(ALU_r_2_), .Q(_601_) );
NO2X1 NO2X1_6 ( .gnd!(gnd!), .vdd!(vdd!), .A(extR[2]), .B(_595__bF_buf0), .Q(_602_) );
ON31X1 ON31X1_3 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_cyc_bF_buf9_bF_buf1), .B(_601_), .C(_602_), .D(_600_), .Q(_6__2_) );
NA2X1 NA2X1_4 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_cyc_bF_buf8_bF_buf0), .B(R_3_), .Q(_603_) );
NO2X1 NO2X1_7 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_IDEC1_cu_custom_inst_bF_buf4), .B(ALU_r_3_), .Q(_604_) );
NO2X1 NO2X1_8 ( .gnd!(gnd!), .vdd!(vdd!), .A(extR[3]), .B(_595__bF_buf0), .Q(_605_) );
ON31X1 ON31X1_4 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_cyc_bF_buf7_bF_buf3), .B(_604_), .C(_605_), .D(_603_), .Q(_6__3_) );
NA2X1 NA2X1_5 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_cyc_bF_buf6_bF_buf0), .B(R_4_), .Q(_606_) );
NO2X1 NO2X1_9 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_IDEC1_cu_custom_inst_bF_buf0), .B(ALU_r_4_), .Q(_607_) );
NO2X1 NO2X1_10 ( .gnd!(gnd!), .vdd!(vdd!), .A(extR[4]), .B(_595__bF_buf3), .Q(_608_) );
ON31X1 ON31X1_5 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_cyc_bF_buf5_bF_buf2), .B(_607_), .C(_608_), .D(_606_), .Q(_6__4_) );
NA2X1 NA2X1_6 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_cyc_bF_buf4_bF_buf0), .B(R_5_), .Q(_609_) );
NO2X1 NO2X1_11 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_IDEC1_cu_custom_inst_bF_buf1), .B(ALU_r_5_), .Q(_610_) );
NO2X1 NO2X1_12 ( .gnd!(gnd!), .vdd!(vdd!), .A(extR[5]), .B(_595__bF_buf0), .Q(_611_) );
ON31X1 ON31X1_6 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_cyc_bF_buf3_bF_buf3), .B(_610_), .C(_611_), .D(_609_), .Q(_6__5_) );
NA2X1 NA2X1_7 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_cyc_bF_buf2_bF_buf2), .B(R_6_), .Q(_612_) );
NO2X1 NO2X1_13 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_IDEC1_cu_custom_inst_bF_buf5), .B(ALU_r_6_), .Q(_613_) );
NO2X1 NO2X1_14 ( .gnd!(gnd!), .vdd!(vdd!), .A(extR[6]), .B(_595__bF_buf2), .Q(_614_) );
ON31X1 ON31X1_7 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_cyc_bF_buf1_bF_buf0), .B(_613_), .C(_614_), .D(_612_), .Q(_6__6_) );
NA2X1 NA2X1_8 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_cyc_bF_buf0_bF_buf3), .B(R_7_), .Q(_615_) );
NO2X1 NO2X1_15 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_IDEC1_cu_custom_inst_bF_buf3), .B(ALU_r_7_), .Q(_616_) );
NO2X1 NO2X1_16 ( .gnd!(gnd!), .vdd!(vdd!), .A(extR[7]), .B(_595__bF_buf1), .Q(_617_) );
ON31X1 ON31X1_8 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_cyc_bF_buf14_bF_buf0), .B(_616_), .C(_617_), .D(_615_), .Q(_6__7_) );
NA2X1 NA2X1_9 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_cyc_bF_buf13_bF_buf0), .B(R_8_), .Q(_618_) );
NO2X1 NO2X1_17 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_IDEC1_cu_custom_inst_bF_buf2), .B(ALU_r_8_), .Q(_619_) );
NO2X1 NO2X1_18 ( .gnd!(gnd!), .vdd!(vdd!), .A(extR[8]), .B(_595__bF_buf3), .Q(_620_) );
ON31X1 ON31X1_9 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_cyc_bF_buf12_bF_buf0), .B(_619_), .C(_620_), .D(_618_), .Q(_6__8_) );
NA2X1 NA2X1_10 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_cyc_bF_buf11_bF_buf0), .B(R_9_), .Q(_621_) );
NO2X1 NO2X1_19 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_IDEC1_cu_custom_inst_bF_buf2), .B(ALU_r_9_), .Q(_622_) );
NO2X1 NO2X1_20 ( .gnd!(gnd!), .vdd!(vdd!), .A(extR[9]), .B(_595__bF_buf3), .Q(_623_) );
ON31X1 ON31X1_10 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_cyc_bF_buf10_bF_buf2), .B(_622_), .C(_623_), .D(_621_), .Q(_6__9_) );
NA2X1 NA2X1_11 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_cyc_bF_buf9_bF_buf0), .B(R_10_), .Q(_624_) );
NO2X1 NO2X1_21 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_IDEC1_cu_custom_inst_bF_buf4), .B(ALU_r_10_), .Q(_625_) );
NO2X1 NO2X1_22 ( .gnd!(gnd!), .vdd!(vdd!), .A(extR[10]), .B(_595__bF_buf0), .Q(_626_) );
ON31X1 ON31X1_11 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_cyc_bF_buf8_bF_buf0), .B(_625_), .C(_626_), .D(_624_), .Q(_6__10_) );
NA2X1 NA2X1_12 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_cyc_bF_buf7_bF_buf1), .B(R_11_), .Q(_627_) );
NO2X1 NO2X1_23 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_IDEC1_cu_custom_inst_bF_buf0), .B(ALU_r_11_), .Q(_628_) );
NO2X1 NO2X1_24 ( .gnd!(gnd!), .vdd!(vdd!), .A(extR[11]), .B(_595__bF_buf3), .Q(_629_) );
ON31X1 ON31X1_12 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_cyc_bF_buf6_bF_buf0), .B(_628_), .C(_629_), .D(_627_), .Q(_6__11_) );
NA2X1 NA2X1_13 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_cyc_bF_buf5_bF_buf2), .B(R_12_), .Q(_630_) );
NO2X1 NO2X1_25 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_IDEC1_cu_custom_inst_bF_buf2), .B(ALU_r_12_), .Q(_631_) );
NO2X1 NO2X1_26 ( .gnd!(gnd!), .vdd!(vdd!), .A(extR[12]), .B(_595__bF_buf2), .Q(_632_) );
ON31X1 ON31X1_13 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_cyc_bF_buf4_bF_buf0), .B(_631_), .C(_632_), .D(_630_), .Q(_6__12_) );
NA2X1 NA2X1_14 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_cyc_bF_buf3_bF_buf3), .B(R_13_), .Q(_633_) );
NO2X1 NO2X1_27 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_IDEC1_cu_custom_inst_bF_buf4), .B(ALU_r_13_), .Q(_634_) );
NO2X1 NO2X1_28 ( .gnd!(gnd!), .vdd!(vdd!), .A(extR[13]), .B(_595__bF_buf1), .Q(_635_) );
ON31X1 ON31X1_14 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_cyc_bF_buf2_bF_buf2), .B(_634_), .C(_635_), .D(_633_), .Q(_6__13_) );
NA2X1 NA2X1_15 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_cyc_bF_buf1_bF_buf0), .B(R_14_), .Q(_636_) );
NO2X1 NO2X1_29 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_IDEC1_cu_custom_inst_bF_buf0), .B(ALU_r_14_), .Q(_637_) );
NO2X1 NO2X1_30 ( .gnd!(gnd!), .vdd!(vdd!), .A(extR[14]), .B(_595__bF_buf2), .Q(_638_) );
ON31X1 ON31X1_15 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_cyc_bF_buf0_bF_buf2), .B(_637_), .C(_638_), .D(_636_), .Q(_6__14_) );
NA2X1 NA2X1_16 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_cyc_bF_buf14_bF_buf0), .B(R_15_), .Q(_639_) );
NO2X1 NO2X1_31 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_IDEC1_cu_custom_inst_bF_buf2), .B(ALU_r_15_), .Q(_640_) );
NO2X1 NO2X1_32 ( .gnd!(gnd!), .vdd!(vdd!), .A(extR[15]), .B(_595__bF_buf1), .Q(_641_) );
ON31X1 ON31X1_16 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_cyc_bF_buf13_bF_buf1), .B(_640_), .C(_641_), .D(_639_), .Q(_6__15_) );
NA2X1 NA2X1_17 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_cyc_bF_buf12_bF_buf3), .B(R_16_), .Q(_642_) );
NO2X1 NO2X1_33 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_IDEC1_cu_custom_inst_bF_buf3), .B(ALU_r_16_), .Q(_643_) );
NO2X1 NO2X1_34 ( .gnd!(gnd!), .vdd!(vdd!), .A(extR[16]), .B(_595__bF_buf4), .Q(_644_) );
ON31X1 ON31X1_17 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_cyc_bF_buf11_bF_buf1), .B(_643_), .C(_644_), .D(_642_), .Q(_6__16_) );
NA2X1 NA2X1_18 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_cyc_bF_buf10_bF_buf2), .B(R_17_), .Q(_645_) );
NO2X1 NO2X1_35 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_IDEC1_cu_custom_inst_bF_buf0), .B(ALU_r_17_), .Q(_646_) );
NO2X1 NO2X1_36 ( .gnd!(gnd!), .vdd!(vdd!), .A(extR[17]), .B(_595__bF_buf3), .Q(_647_) );
ON31X1 ON31X1_18 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_cyc_bF_buf9_bF_buf1), .B(_646_), .C(_647_), .D(_645_), .Q(_6__17_) );
NA2X1 NA2X1_19 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_cyc_bF_buf8_bF_buf2), .B(R_18_), .Q(_648_) );
NO2X1 NO2X1_37 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_IDEC1_cu_custom_inst_bF_buf0), .B(ALU_r_18_), .Q(_649_) );
NO2X1 NO2X1_38 ( .gnd!(gnd!), .vdd!(vdd!), .A(extR[18]), .B(_595__bF_buf3), .Q(_650_) );
ON31X1 ON31X1_19 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_cyc_bF_buf7_bF_buf1), .B(_649_), .C(_650_), .D(_648_), .Q(_6__18_) );
NA2X1 NA2X1_20 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_cyc_bF_buf6_bF_buf2), .B(R_19_), .Q(_651_) );
NO2X1 NO2X1_39 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_IDEC1_cu_custom_inst_bF_buf4), .B(ALU_r_19_), .Q(_652_) );
NO2X1 NO2X1_40 ( .gnd!(gnd!), .vdd!(vdd!), .A(extR[19]), .B(_595__bF_buf0), .Q(_653_) );
ON31X1 ON31X1_20 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_cyc_bF_buf5_bF_buf3), .B(_652_), .C(_653_), .D(_651_), .Q(_6__19_) );
NA2X1 NA2X1_21 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_cyc_bF_buf4_bF_buf0), .B(R_20_), .Q(_654_) );
NO2X1 NO2X1_41 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_IDEC1_cu_custom_inst_bF_buf2), .B(ALU_r_20_), .Q(_655_) );
NO2X1 NO2X1_42 ( .gnd!(gnd!), .vdd!(vdd!), .A(extR[20]), .B(_595__bF_buf1), .Q(_656_) );
ON31X1 ON31X1_21 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_cyc_bF_buf3_bF_buf3), .B(_655_), .C(_656_), .D(_654_), .Q(_6__20_) );
NA2X1 NA2X1_22 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_cyc_bF_buf2_bF_buf2), .B(R_21_), .Q(_657_) );
NO2X1 NO2X1_43 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_IDEC1_cu_custom_inst_bF_buf1), .B(ALU_r_21_), .Q(_658_) );
NO2X1 NO2X1_44 ( .gnd!(gnd!), .vdd!(vdd!), .A(extR[21]), .B(_595__bF_buf4), .Q(_659_) );
ON31X1 ON31X1_22 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_cyc_bF_buf1_bF_buf3), .B(_658_), .C(_659_), .D(_657_), .Q(_6__21_) );
NA2X1 NA2X1_23 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_cyc_bF_buf0_bF_buf3), .B(R_22_), .Q(_660_) );
NO2X1 NO2X1_45 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_IDEC1_cu_custom_inst_bF_buf1), .B(ALU_r_22_), .Q(_661_) );
NO2X1 NO2X1_46 ( .gnd!(gnd!), .vdd!(vdd!), .A(extR[22]), .B(_595__bF_buf4), .Q(_662_) );
ON31X1 ON31X1_23 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_cyc_bF_buf14_bF_buf1), .B(_661_), .C(_662_), .D(_660_), .Q(_6__22_) );
NA2X1 NA2X1_24 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_cyc_bF_buf13_bF_buf2), .B(R_23_), .Q(_663_) );
NO2X1 NO2X1_47 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_IDEC1_cu_custom_inst_bF_buf1), .B(ALU_r_23_), .Q(_664_) );
NO2X1 NO2X1_48 ( .gnd!(gnd!), .vdd!(vdd!), .A(extR[23]), .B(_595__bF_buf4), .Q(_665_) );
ON31X1 ON31X1_24 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_cyc_bF_buf12_bF_buf2), .B(_664_), .C(_665_), .D(_663_), .Q(_6__23_) );
NA2X1 NA2X1_25 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_cyc_bF_buf11_bF_buf0), .B(R_24_), .Q(_666_) );
NO2X1 NO2X1_49 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_IDEC1_cu_custom_inst_bF_buf4), .B(ALU_r_24_), .Q(_667_) );
NO2X1 NO2X1_50 ( .gnd!(gnd!), .vdd!(vdd!), .A(extR[24]), .B(_595__bF_buf3), .Q(_668_) );
ON31X1 ON31X1_25 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_cyc_bF_buf10_bF_buf3), .B(_667_), .C(_668_), .D(_666_), .Q(_6__24_) );
NA2X1 NA2X1_26 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_cyc_bF_buf9_bF_buf1), .B(R_25_), .Q(_669_) );
NO2X1 NO2X1_51 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_IDEC1_cu_custom_inst_bF_buf3), .B(ALU_r_25_), .Q(_670_) );
NO2X1 NO2X1_52 ( .gnd!(gnd!), .vdd!(vdd!), .A(extR[25]), .B(_595__bF_buf4), .Q(_671_) );
ON31X1 ON31X1_26 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_cyc_bF_buf8_bF_buf3), .B(_670_), .C(_671_), .D(_669_), .Q(_6__25_) );
NA2X1 NA2X1_27 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_cyc_bF_buf7_bF_buf3), .B(R_26_), .Q(_672_) );
NO2X1 NO2X1_53 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_IDEC1_cu_custom_inst_bF_buf5), .B(ALU_r_26_), .Q(_673_) );
NO2X1 NO2X1_54 ( .gnd!(gnd!), .vdd!(vdd!), .A(extR[26]), .B(_595__bF_buf1), .Q(_674_) );
ON31X1 ON31X1_27 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_cyc_bF_buf6_bF_buf1), .B(_673_), .C(_674_), .D(_672_), .Q(_6__26_) );
NA2X1 NA2X1_28 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_cyc_bF_buf5_bF_buf1), .B(R_27_), .Q(_675_) );
NO2X1 NO2X1_55 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_IDEC1_cu_custom_inst_bF_buf1), .B(ALU_r_27_), .Q(_676_) );
NO2X1 NO2X1_56 ( .gnd!(gnd!), .vdd!(vdd!), .A(extR[27]), .B(_595__bF_buf4), .Q(_7_) );
ON31X1 ON31X1_28 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_cyc_bF_buf4_bF_buf3), .B(_676_), .C(_7_), .D(_675_), .Q(_6__27_) );
NA2X1 NA2X1_29 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_cyc_bF_buf3_bF_buf2), .B(R_28_), .Q(_8_) );
NO2X1 NO2X1_57 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_IDEC1_cu_custom_inst_bF_buf4), .B(ALU_r_28_), .Q(_9_) );
NO2X1 NO2X1_58 ( .gnd!(gnd!), .vdd!(vdd!), .A(extR[28]), .B(_595__bF_buf0), .Q(_10_) );
ON31X1 ON31X1_29 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_cyc_bF_buf2_bF_buf2), .B(_9_), .C(_10_), .D(_8_), .Q(_6__28_) );
NA2X1 NA2X1_30 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_cyc_bF_buf1_bF_buf0), .B(R_29_), .Q(_11_) );
NO2X1 NO2X1_59 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_IDEC1_cu_custom_inst_bF_buf5), .B(ALU_r_29_), .Q(_12_) );
NO2X1 NO2X1_60 ( .gnd!(gnd!), .vdd!(vdd!), .A(extR[29]), .B(_595__bF_buf2), .Q(_13_) );
ON31X1 ON31X1_30 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_cyc_bF_buf0_bF_buf2), .B(_12_), .C(_13_), .D(_11_), .Q(_6__29_) );
NA2X1 NA2X1_31 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_cyc_bF_buf14_bF_buf3), .B(R_30_), .Q(_14_) );
NO2X1 NO2X1_61 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_IDEC1_cu_custom_inst_bF_buf1), .B(ALU_r_30_), .Q(_15_) );
NO2X1 NO2X1_62 ( .gnd!(gnd!), .vdd!(vdd!), .A(extR[30]), .B(_595__bF_buf4), .Q(_16_) );
ON31X1 ON31X1_31 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_cyc_bF_buf13_bF_buf2), .B(_15_), .C(_16_), .D(_14_), .Q(_6__30_) );
NA2X1 NA2X1_32 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_cyc_bF_buf12_bF_buf1), .B(R_31_), .Q(_17_) );
NO2X1 NO2X1_63 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_IDEC1_cu_custom_inst_bF_buf5), .B(ALU_r_31_), .Q(_18_) );
NO2X1 NO2X1_64 ( .gnd!(gnd!), .vdd!(vdd!), .A(extR[31]), .B(_595__bF_buf1), .Q(_19_) );
ON31X1 ON31X1_32 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_cyc_bF_buf11_bF_buf2), .B(_18_), .C(_19_), .D(_17_), .Q(_6__31_) );
INX1 INX1_1 ( .gnd!(gnd!), .vdd!(vdd!), .A(_678__0_), .Q(_20_) );
INX3 INX3_1 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_cu_r2_ld), .Q(_21_) );
NA2X1 NA2X1_33 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_IDEC1_cu_load_inst_bF_buf4), .B(bdo[0]), .Q(_22_) );
INX3 INX3_2 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_cu_j_inst_1), .Q(_23_) );
NA2I1X1 NA2I1X1_1 ( .gnd!(gnd!), .vdd!(vdd!), .AN(CTRL_IDEC1_cu_system_inst_bF_buf3), .B(R_0_), .Q(_24_) );
NO2I1X1 NO2I1X1_1 ( .gnd!(gnd!), .vdd!(vdd!), .AN(CTRL_cu_csr_rd_s1_bF_buf2), .B(CNTR_Timer_0_), .Q(_25_) );
ON21X1 ON21X1_1 ( .gnd!(gnd!), .vdd!(vdd!), .A(CNTR_Cycle_0_), .B(CTRL_cu_csr_rd_s1_bF_buf2), .C(CTRL_IDEC1_cu_system_inst_bF_buf4), .Q(_26_) );
ON21X1 ON21X1_2 ( .gnd!(gnd!), .vdd!(vdd!), .A(_25_), .B(_26_), .C(_24_), .Q(_27_) );
INX1 INX1_2 ( .gnd!(gnd!), .vdd!(vdd!), .A(PC_0_), .Q(_28_) );
INX3 INX3_3 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_IDEC1_cu_lui_inst), .Q(_29_) );
ON21X1 ON21X1_3 ( .gnd!(gnd!), .vdd!(vdd!), .A(_28_), .B(_23__bF_buf3), .C(_29__bF_buf6), .Q(_30_) );
AN21X1 AN21X1_1 ( .gnd!(gnd!), .vdd!(vdd!), .A(_27_), .B(_23__bF_buf3), .C(_30_), .Q(_31_) );
INX2 INX2_2 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_IDEC1_cu_load_inst_bF_buf1), .Q(_32_) );
ON21X1 ON21X1_4 ( .gnd!(gnd!), .vdd!(vdd!), .A(_29__bF_buf4), .B(I1_0_), .C(_32__bF_buf0), .Q(_33_) );
ON21X1 ON21X1_5 ( .gnd!(gnd!), .vdd!(vdd!), .A(_31_), .B(_33_), .C(_22_), .Q(_34_) );
NA2X1 NA2X1_34 ( .gnd!(gnd!), .vdd!(vdd!), .A(_34_), .B(CTRL_cu_r2_src_bF_buf3), .Q(_35_) );
INX2 INX2_3 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_cu_r2_src_bF_buf1), .Q(_36_) );
NO2X1 NO2X1_65 ( .gnd!(gnd!), .vdd!(vdd!), .A(_687__1_), .B(_687__0_), .Q(_37_) );
NO2X1 NO2X1_66 ( .gnd!(gnd!), .vdd!(vdd!), .A(_687__3_), .B(_687__2_), .Q(_38_) );
NA3I1X2 NA3I1X2_1 ( .gnd!(gnd!), .vdd!(vdd!), .AN(_687__4_), .B(_37_), .C(_38_), .Q(_39_) );
AN31X1 AN31X1_1 ( .gnd!(gnd!), .vdd!(vdd!), .A(_36__bF_buf1), .B(rfRS2[0]), .C(_39__bF_buf3), .D(_21__bF_buf4), .Q(_40_) );
AN22X1 AN22X1_1 ( .gnd!(gnd!), .vdd!(vdd!), .A(_20_), .B(_21__bF_buf4), .C(_35_), .D(_40_), .Q(_4__0_) );
NA2X1 NA2X1_35 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_IDEC1_cu_load_inst_bF_buf0), .B(bdo[1]), .Q(_41_) );
NA2I1X1 NA2I1X1_2 ( .gnd!(gnd!), .vdd!(vdd!), .AN(CTRL_IDEC1_cu_system_inst_bF_buf0), .B(R_1_), .Q(_42_) );
NO2I1X1 NO2I1X1_2 ( .gnd!(gnd!), .vdd!(vdd!), .AN(CTRL_cu_csr_rd_s1_bF_buf2), .B(CNTR_Timer_1_), .Q(_43_) );
ON21X1 ON21X1_6 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_cu_csr_rd_s1_bF_buf5), .B(CNTR_Cycle_1_), .C(CTRL_IDEC1_cu_system_inst_bF_buf1), .Q(_44_) );
ON211X1 ON211X1_1 ( .gnd!(gnd!), .vdd!(vdd!), .A(_43_), .B(_44_), .C(_23__bF_buf6), .D(_42_), .Q(_45_) );
INX1 INX1_3 ( .gnd!(gnd!), .vdd!(vdd!), .A(PC_1_), .Q(_46_) );
NA2X1 NA2X1_36 ( .gnd!(gnd!), .vdd!(vdd!), .A(_46_), .B(CTRL_cu_j_inst_1), .Q(_47_) );
AN21X1 AN21X1_2 ( .gnd!(gnd!), .vdd!(vdd!), .A(_45_), .B(_47_), .C(CTRL_IDEC1_cu_lui_inst), .Q(_48_) );
ON21X1 ON21X1_7 ( .gnd!(gnd!), .vdd!(vdd!), .A(_29__bF_buf0), .B(I1_1_), .C(_32__bF_buf3), .Q(_49_) );
ON211X1 ON211X1_2 ( .gnd!(gnd!), .vdd!(vdd!), .A(_48_), .B(_49_), .C(CTRL_cu_r2_src_bF_buf2), .D(_41_), .Q(_50_) );
AN21X1 AN21X1_3 ( .gnd!(gnd!), .vdd!(vdd!), .A(_39__bF_buf2), .B(rfRS2[1]), .C(CTRL_cu_r2_src_bF_buf3), .Q(_51_) );
NO2X1 NO2X1_67 ( .gnd!(gnd!), .vdd!(vdd!), .A(_21__bF_buf2), .B(_51_), .Q(_52_) );
AO22X2 AO22X2_1 ( .gnd!(gnd!), .vdd!(vdd!), .A(_21__bF_buf6), .B(_678__1_), .C(_50_), .D(_52_), .Q(_4__1_) );
INX1 INX1_4 ( .gnd!(gnd!), .vdd!(vdd!), .A(_678__2_), .Q(_53_) );
NA2X1 NA2X1_37 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_IDEC1_cu_load_inst_bF_buf2), .B(bdo[2]), .Q(_54_) );
NA2I1X1 NA2I1X1_3 ( .gnd!(gnd!), .vdd!(vdd!), .AN(CTRL_IDEC1_cu_system_inst_bF_buf7), .B(R_2_), .Q(_55_) );
NO2I1X1 NO2I1X1_3 ( .gnd!(gnd!), .vdd!(vdd!), .AN(CTRL_cu_csr_rd_s1_bF_buf0), .B(CNTR_Timer_2_), .Q(_56_) );
ON21X1 ON21X1_8 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_cu_csr_rd_s1_bF_buf5), .B(CNTR_Cycle_2_), .C(CTRL_IDEC1_cu_system_inst_bF_buf6), .Q(_57_) );
ON21X1 ON21X1_9 ( .gnd!(gnd!), .vdd!(vdd!), .A(_56_), .B(_57_), .C(_55_), .Q(_58_) );
INX1 INX1_5 ( .gnd!(gnd!), .vdd!(vdd!), .A(PC_2_), .Q(_59_) );
ON21X1 ON21X1_10 ( .gnd!(gnd!), .vdd!(vdd!), .A(_23__bF_buf3), .B(_59_), .C(_29__bF_buf4), .Q(_60_) );
AN21X1 AN21X1_4 ( .gnd!(gnd!), .vdd!(vdd!), .A(_58_), .B(_23__bF_buf1), .C(_60_), .Q(_61_) );
ON21X1 ON21X1_11 ( .gnd!(gnd!), .vdd!(vdd!), .A(_29__bF_buf1), .B(I1_2_), .C(_32__bF_buf2), .Q(_62_) );
ON21X1 ON21X1_12 ( .gnd!(gnd!), .vdd!(vdd!), .A(_61_), .B(_62_), .C(_54_), .Q(_63_) );
NA2X1 NA2X1_38 ( .gnd!(gnd!), .vdd!(vdd!), .A(_63_), .B(CTRL_cu_r2_src_bF_buf3), .Q(_64_) );
AN31X1 AN31X1_2 ( .gnd!(gnd!), .vdd!(vdd!), .A(_36__bF_buf1), .B(rfRS2[2]), .C(_39__bF_buf3), .D(_21__bF_buf4), .Q(_65_) );
AN22X1 AN22X1_2 ( .gnd!(gnd!), .vdd!(vdd!), .A(_21__bF_buf5), .B(_53_), .C(_64_), .D(_65_), .Q(_4__2_) );
NA2X1 NA2X1_39 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_IDEC1_cu_load_inst_bF_buf1), .B(bdo[3]), .Q(_66_) );
NA2I1X1 NA2I1X1_4 ( .gnd!(gnd!), .vdd!(vdd!), .AN(CTRL_IDEC1_cu_system_inst_bF_buf6), .B(R_3_), .Q(_67_) );
NO2I1X1 NO2I1X1_4 ( .gnd!(gnd!), .vdd!(vdd!), .AN(CTRL_cu_csr_rd_s1_bF_buf0), .B(CNTR_Timer_3_), .Q(_68_) );
ON21X1 ON21X1_13 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_cu_csr_rd_s1_bF_buf5), .B(CNTR_Cycle_3_), .C(CTRL_IDEC1_cu_system_inst_bF_buf6), .Q(_69_) );
ON211X1 ON211X1_3 ( .gnd!(gnd!), .vdd!(vdd!), .A(_68_), .B(_69_), .C(_23__bF_buf0), .D(_67_), .Q(_70_) );
INX1 INX1_6 ( .gnd!(gnd!), .vdd!(vdd!), .A(PC_3_), .Q(_71_) );
NA2X1 NA2X1_40 ( .gnd!(gnd!), .vdd!(vdd!), .A(_71_), .B(CTRL_cu_j_inst_1), .Q(_72_) );
AN21X1 AN21X1_5 ( .gnd!(gnd!), .vdd!(vdd!), .A(_70_), .B(_72_), .C(CTRL_IDEC1_cu_lui_inst), .Q(_73_) );
ON21X1 ON21X1_14 ( .gnd!(gnd!), .vdd!(vdd!), .A(_29__bF_buf0), .B(I1_3_), .C(_32__bF_buf3), .Q(_74_) );
ON211X1 ON211X1_4 ( .gnd!(gnd!), .vdd!(vdd!), .A(_73_), .B(_74_), .C(CTRL_cu_r2_src_bF_buf2), .D(_66_), .Q(_75_) );
AN21X1 AN21X1_6 ( .gnd!(gnd!), .vdd!(vdd!), .A(_39__bF_buf3), .B(rfRS2[3]), .C(CTRL_cu_r2_src_bF_buf3), .Q(_76_) );
NO2X1 NO2X1_68 ( .gnd!(gnd!), .vdd!(vdd!), .A(_21__bF_buf5), .B(_76_), .Q(_77_) );
AO22X2 AO22X2_2 ( .gnd!(gnd!), .vdd!(vdd!), .A(_21__bF_buf5), .B(_678__3_), .C(_75_), .D(_77_), .Q(_4__3_) );
INX1 INX1_7 ( .gnd!(gnd!), .vdd!(vdd!), .A(_678__4_), .Q(_78_) );
NA2X1 NA2X1_41 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_IDEC1_cu_load_inst_bF_buf3), .B(bdo[4]), .Q(_79_) );
NA2I1X1 NA2I1X1_5 ( .gnd!(gnd!), .vdd!(vdd!), .AN(CTRL_IDEC1_cu_system_inst_bF_buf4), .B(R_4_), .Q(_80_) );
NO2I1X1 NO2I1X1_5 ( .gnd!(gnd!), .vdd!(vdd!), .AN(CTRL_cu_csr_rd_s1_bF_buf0), .B(CNTR_Timer_4_), .Q(_81_) );
ON21X1 ON21X1_15 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_cu_csr_rd_s1_bF_buf0), .B(CNTR_Cycle_4_), .C(CTRL_IDEC1_cu_system_inst_bF_buf4), .Q(_82_) );
ON21X1 ON21X1_16 ( .gnd!(gnd!), .vdd!(vdd!), .A(_81_), .B(_82_), .C(_80_), .Q(_83_) );
INX1 INX1_8 ( .gnd!(gnd!), .vdd!(vdd!), .A(PC_4_), .Q(_84_) );
ON21X1 ON21X1_17 ( .gnd!(gnd!), .vdd!(vdd!), .A(_23__bF_buf1), .B(_84_), .C(_29__bF_buf2), .Q(_85_) );
AN21X1 AN21X1_7 ( .gnd!(gnd!), .vdd!(vdd!), .A(_83_), .B(_23__bF_buf1), .C(_85_), .Q(_86_) );
ON21X1 ON21X1_18 ( .gnd!(gnd!), .vdd!(vdd!), .A(_29__bF_buf4), .B(I1_4_), .C(_32__bF_buf0), .Q(_87_) );
ON21X1 ON21X1_19 ( .gnd!(gnd!), .vdd!(vdd!), .A(_86_), .B(_87_), .C(_79_), .Q(_88_) );
NA2X1 NA2X1_42 ( .gnd!(gnd!), .vdd!(vdd!), .A(_88_), .B(CTRL_cu_r2_src_bF_buf0), .Q(_89_) );
AN31X1 AN31X1_3 ( .gnd!(gnd!), .vdd!(vdd!), .A(_36__bF_buf2), .B(rfRS2[4]), .C(_39__bF_buf4), .D(_21__bF_buf1), .Q(_90_) );
AN22X1 AN22X1_3 ( .gnd!(gnd!), .vdd!(vdd!), .A(_21__bF_buf1), .B(_78_), .C(_89_), .D(_90_), .Q(_4__4_) );
NA2X1 NA2X1_43 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_IDEC1_cu_load_inst_bF_buf1), .B(bdo[5]), .Q(_91_) );
NA2I1X1 NA2I1X1_6 ( .gnd!(gnd!), .vdd!(vdd!), .AN(CTRL_IDEC1_cu_system_inst_bF_buf4), .B(R_5_), .Q(_92_) );
NO2I1X1 NO2I1X1_6 ( .gnd!(gnd!), .vdd!(vdd!), .AN(CTRL_cu_csr_rd_s1_bF_buf1), .B(CNTR_Timer_5_), .Q(_93_) );
ON21X1 ON21X1_20 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_cu_csr_rd_s1_bF_buf1), .B(CNTR_Cycle_5_), .C(CTRL_IDEC1_cu_system_inst_bF_buf5), .Q(_94_) );
ON211X1 ON211X1_5 ( .gnd!(gnd!), .vdd!(vdd!), .A(_93_), .B(_94_), .C(_23__bF_buf4), .D(_92_), .Q(_95_) );
INX1 INX1_9 ( .gnd!(gnd!), .vdd!(vdd!), .A(PC_5_), .Q(_96_) );
NA2X1 NA2X1_44 ( .gnd!(gnd!), .vdd!(vdd!), .A(_96_), .B(CTRL_cu_j_inst_1), .Q(_97_) );
AN21X1 AN21X1_8 ( .gnd!(gnd!), .vdd!(vdd!), .A(_95_), .B(_97_), .C(CTRL_IDEC1_cu_lui_inst), .Q(_98_) );
ON21X1 ON21X1_21 ( .gnd!(gnd!), .vdd!(vdd!), .A(_29__bF_buf0), .B(I1_5_), .C(_32__bF_buf3), .Q(_99_) );
ON211X1 ON211X1_6 ( .gnd!(gnd!), .vdd!(vdd!), .A(_98_), .B(_99_), .C(CTRL_cu_r2_src_bF_buf2), .D(_91_), .Q(_100_) );
AN21X1 AN21X1_9 ( .gnd!(gnd!), .vdd!(vdd!), .A(_39__bF_buf0), .B(rfRS2[5]), .C(CTRL_cu_r2_src_bF_buf1), .Q(_101_) );
NO2X1 NO2X1_69 ( .gnd!(gnd!), .vdd!(vdd!), .A(_21__bF_buf2), .B(_101_), .Q(_102_) );
AO22X2 AO22X2_3 ( .gnd!(gnd!), .vdd!(vdd!), .A(_21__bF_buf6), .B(_678__5_), .C(_100_), .D(_102_), .Q(_4__5_) );
INX1 INX1_10 ( .gnd!(gnd!), .vdd!(vdd!), .A(_678__6_), .Q(_103_) );
NA2X1 NA2X1_45 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_IDEC1_cu_load_inst_bF_buf4), .B(bdo[6]), .Q(_104_) );
NA2I1X1 NA2I1X1_7 ( .gnd!(gnd!), .vdd!(vdd!), .AN(CTRL_IDEC1_cu_system_inst_bF_buf3), .B(R_6_), .Q(_105_) );
NO2I1X1 NO2I1X1_7 ( .gnd!(gnd!), .vdd!(vdd!), .AN(CTRL_cu_csr_rd_s1_bF_buf0), .B(CNTR_Timer_6_), .Q(_106_) );
ON21X1 ON21X1_22 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_cu_csr_rd_s1_bF_buf0), .B(CNTR_Cycle_6_), .C(CTRL_IDEC1_cu_system_inst_bF_buf4), .Q(_107_) );
ON21X1 ON21X1_23 ( .gnd!(gnd!), .vdd!(vdd!), .A(_106_), .B(_107_), .C(_105_), .Q(_108_) );
INX1 INX1_11 ( .gnd!(gnd!), .vdd!(vdd!), .A(PC_6_), .Q(_109_) );
ON21X1 ON21X1_24 ( .gnd!(gnd!), .vdd!(vdd!), .A(_23__bF_buf5), .B(_109_), .C(_29__bF_buf6), .Q(_110_) );
AN21X1 AN21X1_10 ( .gnd!(gnd!), .vdd!(vdd!), .A(_108_), .B(_23__bF_buf5), .C(_110_), .Q(_111_) );
ON21X1 ON21X1_25 ( .gnd!(gnd!), .vdd!(vdd!), .A(_29__bF_buf5), .B(I1_6_), .C(_32__bF_buf2), .Q(_112_) );
ON21X1 ON21X1_26 ( .gnd!(gnd!), .vdd!(vdd!), .A(_111_), .B(_112_), .C(_104_), .Q(_113_) );
NA2X1 NA2X1_46 ( .gnd!(gnd!), .vdd!(vdd!), .A(_113_), .B(CTRL_cu_r2_src_bF_buf2), .Q(_114_) );
AN31X1 AN31X1_4 ( .gnd!(gnd!), .vdd!(vdd!), .A(_36__bF_buf3), .B(rfRS2[6]), .C(_39__bF_buf1), .D(_21__bF_buf3), .Q(_115_) );
AN22X1 AN22X1_4 ( .gnd!(gnd!), .vdd!(vdd!), .A(_21__bF_buf3), .B(_103_), .C(_114_), .D(_115_), .Q(_4__6_) );
NA2X1 NA2X1_47 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_IDEC1_cu_load_inst_bF_buf2), .B(bdo[7]), .Q(_116_) );
NA2I1X1 NA2I1X1_8 ( .gnd!(gnd!), .vdd!(vdd!), .AN(CTRL_IDEC1_cu_system_inst_bF_buf4), .B(R_7_), .Q(_117_) );
NO2I1X1 NO2I1X1_8 ( .gnd!(gnd!), .vdd!(vdd!), .AN(CTRL_cu_csr_rd_s1_bF_buf0), .B(CNTR_Timer_7_), .Q(_118_) );
ON21X1 ON21X1_27 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_cu_csr_rd_s1_bF_buf1), .B(CNTR_Cycle_7_), .C(CTRL_IDEC1_cu_system_inst_bF_buf5), .Q(_119_) );
ON211X1 ON211X1_7 ( .gnd!(gnd!), .vdd!(vdd!), .A(_118_), .B(_119_), .C(_23__bF_buf4), .D(_117_), .Q(_120_) );
INX1 INX1_12 ( .gnd!(gnd!), .vdd!(vdd!), .A(PC_7_), .Q(_121_) );
NA2X1 NA2X1_48 ( .gnd!(gnd!), .vdd!(vdd!), .A(_121_), .B(CTRL_cu_j_inst_1), .Q(_122_) );
AN21X1 AN21X1_11 ( .gnd!(gnd!), .vdd!(vdd!), .A(_120_), .B(_122_), .C(CTRL_IDEC1_cu_lui_inst), .Q(_123_) );
ON21X1 ON21X1_28 ( .gnd!(gnd!), .vdd!(vdd!), .A(_29__bF_buf1), .B(I1_7_), .C(_32__bF_buf1), .Q(_124_) );
ON211X1 ON211X1_8 ( .gnd!(gnd!), .vdd!(vdd!), .A(_123_), .B(_124_), .C(CTRL_cu_r2_src_bF_buf5), .D(_116_), .Q(_125_) );
NA2X1 NA2X1_49 ( .gnd!(gnd!), .vdd!(vdd!), .A(_39__bF_buf0), .B(rfRS2[7]), .Q(_126_) );
AN21X1 AN21X1_12 ( .gnd!(gnd!), .vdd!(vdd!), .A(_126_), .B(_36__bF_buf0), .C(_21__bF_buf1), .Q(_127_) );
AO22X2 AO22X2_4 ( .gnd!(gnd!), .vdd!(vdd!), .A(_21__bF_buf2), .B(_678__7_), .C(_125_), .D(_127_), .Q(_4__7_) );
NA2X1 NA2X1_50 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_IDEC1_cu_load_inst_bF_buf1), .B(EXT_do_8_), .Q(_128_) );
NA2I1X1 NA2I1X1_9 ( .gnd!(gnd!), .vdd!(vdd!), .AN(CTRL_IDEC1_cu_system_inst_bF_buf0), .B(R_8_), .Q(_129_) );
NO2I1X1 NO2I1X1_9 ( .gnd!(gnd!), .vdd!(vdd!), .AN(CTRL_cu_csr_rd_s1_bF_buf7), .B(CNTR_Timer_8_), .Q(_130_) );
ON21X1 ON21X1_29 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_cu_csr_rd_s1_bF_buf6), .B(CNTR_Cycle_8_), .C(CTRL_IDEC1_cu_system_inst_bF_buf1), .Q(_131_) );
ON211X1 ON211X1_9 ( .gnd!(gnd!), .vdd!(vdd!), .A(_130_), .B(_131_), .C(_23__bF_buf0), .D(_129_), .Q(_132_) );
INX1 INX1_13 ( .gnd!(gnd!), .vdd!(vdd!), .A(PC_8_), .Q(_133_) );
NA2X1 NA2X1_51 ( .gnd!(gnd!), .vdd!(vdd!), .A(_133_), .B(CTRL_cu_j_inst_1), .Q(_134_) );
AN21X1 AN21X1_13 ( .gnd!(gnd!), .vdd!(vdd!), .A(_132_), .B(_134_), .C(CTRL_IDEC1_cu_lui_inst), .Q(_135_) );
ON21X1 ON21X1_30 ( .gnd!(gnd!), .vdd!(vdd!), .A(_29__bF_buf0), .B(I1_8_), .C(_32__bF_buf3), .Q(_136_) );
ON211X1 ON211X1_10 ( .gnd!(gnd!), .vdd!(vdd!), .A(_135_), .B(_136_), .C(CTRL_cu_r2_src_bF_buf5), .D(_128_), .Q(_137_) );
AN21X1 AN21X1_14 ( .gnd!(gnd!), .vdd!(vdd!), .A(_39__bF_buf3), .B(rfRS2[8]), .C(CTRL_cu_r2_src_bF_buf3), .Q(_138_) );
NO2X1 NO2X1_70 ( .gnd!(gnd!), .vdd!(vdd!), .A(_21__bF_buf5), .B(_138_), .Q(_139_) );
AO22X2 AO22X2_5 ( .gnd!(gnd!), .vdd!(vdd!), .A(_21__bF_buf2), .B(_678__8_), .C(_137_), .D(_139_), .Q(_4__8_) );
INX1 INX1_14 ( .gnd!(gnd!), .vdd!(vdd!), .A(_678__9_), .Q(_140_) );
NA2X1 NA2X1_52 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_IDEC1_cu_load_inst_bF_buf0), .B(EXT_do_9_), .Q(_141_) );
NA2I1X1 NA2I1X1_10 ( .gnd!(gnd!), .vdd!(vdd!), .AN(CTRL_IDEC1_cu_system_inst_bF_buf7), .B(R_9_), .Q(_142_) );
NO2I1X1 NO2I1X1_10 ( .gnd!(gnd!), .vdd!(vdd!), .AN(CTRL_cu_csr_rd_s1_bF_buf1), .B(CNTR_Timer_9_), .Q(_143_) );
ON21X1 ON21X1_31 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_cu_csr_rd_s1_bF_buf3), .B(CNTR_Cycle_9_), .C(CTRL_IDEC1_cu_system_inst_bF_buf5), .Q(_144_) );
ON21X1 ON21X1_32 ( .gnd!(gnd!), .vdd!(vdd!), .A(_143_), .B(_144_), .C(_142_), .Q(_145_) );
INX1 INX1_15 ( .gnd!(gnd!), .vdd!(vdd!), .A(PC_9_), .Q(_146_) );
ON21X1 ON21X1_33 ( .gnd!(gnd!), .vdd!(vdd!), .A(_23__bF_buf6), .B(_146_), .C(_29__bF_buf5), .Q(_147_) );
AN21X1 AN21X1_15 ( .gnd!(gnd!), .vdd!(vdd!), .A(_145_), .B(_23__bF_buf0), .C(_147_), .Q(_148_) );
ON21X1 ON21X1_34 ( .gnd!(gnd!), .vdd!(vdd!), .A(_29__bF_buf1), .B(I1_9_), .C(_32__bF_buf1), .Q(_149_) );
ON21X1 ON21X1_35 ( .gnd!(gnd!), .vdd!(vdd!), .A(_148_), .B(_149_), .C(_141_), .Q(_150_) );
NA2X1 NA2X1_53 ( .gnd!(gnd!), .vdd!(vdd!), .A(_150_), .B(CTRL_cu_r2_src_bF_buf4), .Q(_151_) );
AN31X1 AN31X1_5 ( .gnd!(gnd!), .vdd!(vdd!), .A(_36__bF_buf0), .B(rfRS2[9]), .C(_39__bF_buf0), .D(_21__bF_buf1), .Q(_152_) );
AN22X1 AN22X1_5 ( .gnd!(gnd!), .vdd!(vdd!), .A(_21__bF_buf2), .B(_140_), .C(_151_), .D(_152_), .Q(_4__9_) );
INX1 INX1_16 ( .gnd!(gnd!), .vdd!(vdd!), .A(_678__10_), .Q(_153_) );
NA2X1 NA2X1_54 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_IDEC1_cu_load_inst_bF_buf3), .B(EXT_do_10_), .Q(_154_) );
NA2I1X1 NA2I1X1_11 ( .gnd!(gnd!), .vdd!(vdd!), .AN(CTRL_IDEC1_cu_system_inst_bF_buf0), .B(R_10_), .Q(_155_) );
NO2I1X1 NO2I1X1_11 ( .gnd!(gnd!), .vdd!(vdd!), .AN(CTRL_cu_csr_rd_s1_bF_buf7), .B(CNTR_Timer_10_), .Q(_156_) );
ON21X1 ON21X1_36 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_cu_csr_rd_s1_bF_buf6), .B(CNTR_Cycle_10_), .C(CTRL_IDEC1_cu_system_inst_bF_buf1), .Q(_157_) );
ON21X1 ON21X1_37 ( .gnd!(gnd!), .vdd!(vdd!), .A(_156_), .B(_157_), .C(_155_), .Q(_158_) );
INX1 INX1_17 ( .gnd!(gnd!), .vdd!(vdd!), .A(PC_10_), .Q(_159_) );
ON21X1 ON21X1_38 ( .gnd!(gnd!), .vdd!(vdd!), .A(_23__bF_buf3), .B(_159_), .C(_29__bF_buf4), .Q(_160_) );
AN21X1 AN21X1_16 ( .gnd!(gnd!), .vdd!(vdd!), .A(_158_), .B(_23__bF_buf0), .C(_160_), .Q(_161_) );
ON21X1 ON21X1_39 ( .gnd!(gnd!), .vdd!(vdd!), .A(_29__bF_buf1), .B(I1_10_), .C(_32__bF_buf1), .Q(_162_) );
ON21X1 ON21X1_40 ( .gnd!(gnd!), .vdd!(vdd!), .A(_161_), .B(_162_), .C(_154_), .Q(_163_) );
NA2X1 NA2X1_55 ( .gnd!(gnd!), .vdd!(vdd!), .A(_163_), .B(CTRL_cu_r2_src_bF_buf1), .Q(_164_) );
AN31X1 AN31X1_6 ( .gnd!(gnd!), .vdd!(vdd!), .A(_36__bF_buf1), .B(rfRS2[10]), .C(_39__bF_buf4), .D(_21__bF_buf4), .Q(_165_) );
AN22X1 AN22X1_6 ( .gnd!(gnd!), .vdd!(vdd!), .A(_21__bF_buf0), .B(_153_), .C(_164_), .D(_165_), .Q(_4__10_) );
INX1 INX1_18 ( .gnd!(gnd!), .vdd!(vdd!), .A(_678__11_), .Q(_166_) );
NA2X1 NA2X1_56 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_IDEC1_cu_load_inst_bF_buf0), .B(EXT_do_11_), .Q(_167_) );
NA2I1X1 NA2I1X1_12 ( .gnd!(gnd!), .vdd!(vdd!), .AN(CTRL_IDEC1_cu_system_inst_bF_buf3), .B(R_11_), .Q(_168_) );
NO2I1X1 NO2I1X1_12 ( .gnd!(gnd!), .vdd!(vdd!), .AN(CTRL_cu_csr_rd_s1_bF_buf4), .B(CNTR_Timer_11_), .Q(_169_) );
ON21X1 ON21X1_41 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_cu_csr_rd_s1_bF_buf3), .B(CNTR_Cycle_11_), .C(CTRL_IDEC1_cu_system_inst_bF_buf5), .Q(_170_) );
ON21X1 ON21X1_42 ( .gnd!(gnd!), .vdd!(vdd!), .A(_169_), .B(_170_), .C(_168_), .Q(_171_) );
INX1 INX1_19 ( .gnd!(gnd!), .vdd!(vdd!), .A(PC_11_), .Q(_172_) );
ON21X1 ON21X1_43 ( .gnd!(gnd!), .vdd!(vdd!), .A(_23__bF_buf1), .B(_172_), .C(_29__bF_buf2), .Q(_173_) );
AN21X1 AN21X1_17 ( .gnd!(gnd!), .vdd!(vdd!), .A(_171_), .B(_23__bF_buf1), .C(_173_), .Q(_174_) );
ON21X1 ON21X1_44 ( .gnd!(gnd!), .vdd!(vdd!), .A(_29__bF_buf5), .B(I1_11_), .C(_32__bF_buf2), .Q(_175_) );
ON21X1 ON21X1_45 ( .gnd!(gnd!), .vdd!(vdd!), .A(_174_), .B(_175_), .C(_167_), .Q(_176_) );
NA2X1 NA2X1_57 ( .gnd!(gnd!), .vdd!(vdd!), .A(_176_), .B(CTRL_cu_r2_src_bF_buf1), .Q(_177_) );
AN31X1 AN31X1_7 ( .gnd!(gnd!), .vdd!(vdd!), .A(_36__bF_buf2), .B(rfRS2[11]), .C(_39__bF_buf4), .D(_21__bF_buf4), .Q(_178_) );
AN22X1 AN22X1_7 ( .gnd!(gnd!), .vdd!(vdd!), .A(_21__bF_buf4), .B(_166_), .C(_177_), .D(_178_), .Q(_4__11_) );
INX1 INX1_20 ( .gnd!(gnd!), .vdd!(vdd!), .A(_678__12_), .Q(_179_) );
NA2X1 NA2X1_58 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_IDEC1_cu_load_inst_bF_buf2), .B(EXT_do_12_), .Q(_180_) );
NA2I1X1 NA2I1X1_13 ( .gnd!(gnd!), .vdd!(vdd!), .AN(CTRL_IDEC1_cu_system_inst_bF_buf3), .B(R_12_), .Q(_181_) );
NO2I1X1 NO2I1X1_13 ( .gnd!(gnd!), .vdd!(vdd!), .AN(CTRL_cu_csr_rd_s1_bF_buf4), .B(CNTR_Timer_12_), .Q(_182_) );
ON21X1 ON21X1_46 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_cu_csr_rd_s1_bF_buf4), .B(CNTR_Cycle_12_), .C(CTRL_IDEC1_cu_system_inst_bF_buf5), .Q(_183_) );
ON21X1 ON21X1_47 ( .gnd!(gnd!), .vdd!(vdd!), .A(_182_), .B(_183_), .C(_181_), .Q(_184_) );
INX1 INX1_21 ( .gnd!(gnd!), .vdd!(vdd!), .A(PC_12_), .Q(_185_) );
ON21X1 ON21X1_48 ( .gnd!(gnd!), .vdd!(vdd!), .A(_23__bF_buf5), .B(_185_), .C(_29__bF_buf2), .Q(_186_) );
AN21X1 AN21X1_18 ( .gnd!(gnd!), .vdd!(vdd!), .A(_184_), .B(_23__bF_buf4), .C(_186_), .Q(_187_) );
ON21X1 ON21X1_49 ( .gnd!(gnd!), .vdd!(vdd!), .A(_29__bF_buf1), .B(I1_12_), .C(_32__bF_buf1), .Q(_188_) );
ON21X1 ON21X1_50 ( .gnd!(gnd!), .vdd!(vdd!), .A(_187_), .B(_188_), .C(_180_), .Q(_189_) );
NA2X1 NA2X1_59 ( .gnd!(gnd!), .vdd!(vdd!), .A(_189_), .B(CTRL_cu_r2_src_bF_buf0), .Q(_190_) );
AN31X1 AN31X1_8 ( .gnd!(gnd!), .vdd!(vdd!), .A(_36__bF_buf2), .B(rfRS2[12]), .C(_39__bF_buf4), .D(_21__bF_buf4), .Q(_191_) );
AN22X1 AN22X1_8 ( .gnd!(gnd!), .vdd!(vdd!), .A(_21__bF_buf0), .B(_179_), .C(_190_), .D(_191_), .Q(_4__12_) );
NA2X1 NA2X1_60 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_IDEC1_cu_load_inst_bF_buf2), .B(EXT_do_13_), .Q(_192_) );
NA2I1X1 NA2I1X1_14 ( .gnd!(gnd!), .vdd!(vdd!), .AN(CTRL_IDEC1_cu_system_inst_bF_buf2), .B(R_13_), .Q(_193_) );
NO2I1X1 NO2I1X1_14 ( .gnd!(gnd!), .vdd!(vdd!), .AN(CTRL_cu_csr_rd_s1_bF_buf3), .B(CNTR_Timer_13_), .Q(_194_) );
ON21X1 ON21X1_51 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_cu_csr_rd_s1_bF_buf3), .B(CNTR_Cycle_13_), .C(CTRL_IDEC1_cu_system_inst_bF_buf2), .Q(_195_) );
ON211X1 ON211X1_11 ( .gnd!(gnd!), .vdd!(vdd!), .A(_194_), .B(_195_), .C(_23__bF_buf4), .D(_193_), .Q(_196_) );
INX1 INX1_22 ( .gnd!(gnd!), .vdd!(vdd!), .A(PC_13_), .Q(_197_) );
NA2X1 NA2X1_61 ( .gnd!(gnd!), .vdd!(vdd!), .A(_197_), .B(CTRL_cu_j_inst_1), .Q(_198_) );
AN21X1 AN21X1_19 ( .gnd!(gnd!), .vdd!(vdd!), .A(_196_), .B(_198_), .C(CTRL_IDEC1_cu_lui_inst), .Q(_199_) );
ON21X1 ON21X1_52 ( .gnd!(gnd!), .vdd!(vdd!), .A(_29__bF_buf0), .B(I1_13_), .C(_32__bF_buf3), .Q(_200_) );
ON211X1 ON211X1_12 ( .gnd!(gnd!), .vdd!(vdd!), .A(_199_), .B(_200_), .C(CTRL_cu_r2_src_bF_buf5), .D(_192_), .Q(_201_) );
AN21X1 AN21X1_20 ( .gnd!(gnd!), .vdd!(vdd!), .A(_39__bF_buf3), .B(rfRS2[13]), .C(CTRL_cu_r2_src_bF_buf3), .Q(_202_) );
NO2X1 NO2X1_71 ( .gnd!(gnd!), .vdd!(vdd!), .A(_21__bF_buf5), .B(_202_), .Q(_203_) );
AO22X2 AO22X2_6 ( .gnd!(gnd!), .vdd!(vdd!), .A(_21__bF_buf2), .B(_678__13_), .C(_201_), .D(_203_), .Q(_4__13_) );
INX1 INX1_23 ( .gnd!(gnd!), .vdd!(vdd!), .A(_678__14_), .Q(_204_) );
NA2X1 NA2X1_62 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_IDEC1_cu_load_inst_bF_buf0), .B(EXT_do_14_), .Q(_205_) );
NA2I1X1 NA2I1X1_15 ( .gnd!(gnd!), .vdd!(vdd!), .AN(CTRL_IDEC1_cu_system_inst_bF_buf7), .B(R_14_), .Q(_206_) );
NO2I1X1 NO2I1X1_15 ( .gnd!(gnd!), .vdd!(vdd!), .AN(CTRL_cu_csr_rd_s1_bF_buf0), .B(CNTR_Timer_14_), .Q(_207_) );
ON21X1 ON21X1_53 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_cu_csr_rd_s1_bF_buf3), .B(CNTR_Cycle_14_), .C(CTRL_IDEC1_cu_system_inst_bF_buf5), .Q(_208_) );
ON21X1 ON21X1_54 ( .gnd!(gnd!), .vdd!(vdd!), .A(_207_), .B(_208_), .C(_206_), .Q(_209_) );
INX1 INX1_24 ( .gnd!(gnd!), .vdd!(vdd!), .A(PC_14_), .Q(_210_) );
ON21X1 ON21X1_55 ( .gnd!(gnd!), .vdd!(vdd!), .A(_23__bF_buf5), .B(_210_), .C(_29__bF_buf2), .Q(_211_) );
AN21X1 AN21X1_21 ( .gnd!(gnd!), .vdd!(vdd!), .A(_209_), .B(_23__bF_buf4), .C(_211_), .Q(_212_) );
ON21X1 ON21X1_56 ( .gnd!(gnd!), .vdd!(vdd!), .A(_29__bF_buf1), .B(I1_14_), .C(_32__bF_buf1), .Q(_213_) );
ON21X1 ON21X1_57 ( .gnd!(gnd!), .vdd!(vdd!), .A(_212_), .B(_213_), .C(_205_), .Q(_214_) );
NA2X1 NA2X1_63 ( .gnd!(gnd!), .vdd!(vdd!), .A(_214_), .B(CTRL_cu_r2_src_bF_buf4), .Q(_215_) );
AN31X1 AN31X1_9 ( .gnd!(gnd!), .vdd!(vdd!), .A(_36__bF_buf1), .B(rfRS2[14]), .C(_39__bF_buf3), .D(_21__bF_buf5), .Q(_216_) );
AN22X1 AN22X1_9 ( .gnd!(gnd!), .vdd!(vdd!), .A(_21__bF_buf5), .B(_204_), .C(_215_), .D(_216_), .Q(_4__14_) );
INX1 INX1_25 ( .gnd!(gnd!), .vdd!(vdd!), .A(_678__15_), .Q(_217_) );
NA2X1 NA2X1_64 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_IDEC1_cu_load_inst_bF_buf3), .B(EXT_do_15_), .Q(_218_) );
NA2I1X1 NA2I1X1_16 ( .gnd!(gnd!), .vdd!(vdd!), .AN(CTRL_IDEC1_cu_system_inst_bF_buf4), .B(R_15_), .Q(_219_) );
NO2I1X1 NO2I1X1_16 ( .gnd!(gnd!), .vdd!(vdd!), .AN(CTRL_cu_csr_rd_s1_bF_buf2), .B(CNTR_Timer_15_), .Q(_220_) );
ON21X1 ON21X1_58 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_cu_csr_rd_s1_bF_buf2), .B(CNTR_Cycle_15_), .C(CTRL_IDEC1_cu_system_inst_bF_buf4), .Q(_221_) );
ON21X1 ON21X1_59 ( .gnd!(gnd!), .vdd!(vdd!), .A(_220_), .B(_221_), .C(_219_), .Q(_222_) );
INX1 INX1_26 ( .gnd!(gnd!), .vdd!(vdd!), .A(PC_15_), .Q(_223_) );
ON21X1 ON21X1_60 ( .gnd!(gnd!), .vdd!(vdd!), .A(_23__bF_buf5), .B(_223_), .C(_29__bF_buf2), .Q(_224_) );
AN21X1 AN21X1_22 ( .gnd!(gnd!), .vdd!(vdd!), .A(_222_), .B(_23__bF_buf5), .C(_224_), .Q(_225_) );
ON21X1 ON21X1_61 ( .gnd!(gnd!), .vdd!(vdd!), .A(_29__bF_buf5), .B(I1_15_), .C(_32__bF_buf2), .Q(_226_) );
ON21X1 ON21X1_62 ( .gnd!(gnd!), .vdd!(vdd!), .A(_225_), .B(_226_), .C(_218_), .Q(_227_) );
NA2X1 NA2X1_65 ( .gnd!(gnd!), .vdd!(vdd!), .A(_227_), .B(CTRL_cu_r2_src_bF_buf4), .Q(_228_) );
AN31X1 AN31X1_10 ( .gnd!(gnd!), .vdd!(vdd!), .A(_36__bF_buf1), .B(rfRS2[15]), .C(_39__bF_buf3), .D(_21__bF_buf4), .Q(_229_) );
AN22X1 AN22X1_10 ( .gnd!(gnd!), .vdd!(vdd!), .A(_21__bF_buf5), .B(_217_), .C(_228_), .D(_229_), .Q(_4__15_) );
NA2X1 NA2X1_66 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_IDEC1_cu_load_inst_bF_buf4), .B(EXT_do_16_), .Q(_230_) );
NA2I1X1 NA2I1X1_17 ( .gnd!(gnd!), .vdd!(vdd!), .AN(CTRL_IDEC1_cu_system_inst_bF_buf6), .B(R_16_), .Q(_231_) );
NO2I1X1 NO2I1X1_17 ( .gnd!(gnd!), .vdd!(vdd!), .AN(CTRL_cu_csr_rd_s1_bF_buf3), .B(CNTR_Timer_16_), .Q(_232_) );
ON21X1 ON21X1_63 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_cu_csr_rd_s1_bF_buf5), .B(CNTR_Cycle_16_), .C(CTRL_IDEC1_cu_system_inst_bF_buf6), .Q(_233_) );
ON211X1 ON211X1_13 ( .gnd!(gnd!), .vdd!(vdd!), .A(_232_), .B(_233_), .C(_23__bF_buf0), .D(_231_), .Q(_234_) );
INX1 INX1_27 ( .gnd!(gnd!), .vdd!(vdd!), .A(PC_16_), .Q(_235_) );
NA2X1 NA2X1_67 ( .gnd!(gnd!), .vdd!(vdd!), .A(_235_), .B(CTRL_cu_j_inst_1), .Q(_236_) );
AN21X1 AN21X1_23 ( .gnd!(gnd!), .vdd!(vdd!), .A(_234_), .B(_236_), .C(CTRL_IDEC1_cu_lui_inst), .Q(_237_) );
ON21X1 ON21X1_64 ( .gnd!(gnd!), .vdd!(vdd!), .A(_29__bF_buf1), .B(I1_16_), .C(_32__bF_buf1), .Q(_238_) );
ON211X1 ON211X1_14 ( .gnd!(gnd!), .vdd!(vdd!), .A(_237_), .B(_238_), .C(CTRL_cu_r2_src_bF_buf5), .D(_230_), .Q(_239_) );
NA2X1 NA2X1_68 ( .gnd!(gnd!), .vdd!(vdd!), .A(_39__bF_buf0), .B(rfRS2[16]), .Q(_240_) );
AN21X1 AN21X1_24 ( .gnd!(gnd!), .vdd!(vdd!), .A(_240_), .B(_36__bF_buf3), .C(_21__bF_buf7), .Q(_241_) );
AO22X2 AO22X2_7 ( .gnd!(gnd!), .vdd!(vdd!), .A(_21__bF_buf3), .B(_678__16_), .C(_239_), .D(_241_), .Q(_4__16_) );
INX1 INX1_28 ( .gnd!(gnd!), .vdd!(vdd!), .A(_678__17_), .Q(_242_) );
NA2X1 NA2X1_69 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_IDEC1_cu_load_inst_bF_buf0), .B(EXT_do_17_), .Q(_243_) );
NA2I1X1 NA2I1X1_18 ( .gnd!(gnd!), .vdd!(vdd!), .AN(CTRL_IDEC1_cu_system_inst_bF_buf7), .B(R_17_), .Q(_244_) );
NO2I1X1 NO2I1X1_18 ( .gnd!(gnd!), .vdd!(vdd!), .AN(CTRL_cu_csr_rd_s1_bF_buf7), .B(CNTR_Timer_17_), .Q(_245_) );
ON21X1 ON21X1_65 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_cu_csr_rd_s1_bF_buf5), .B(CNTR_Cycle_17_), .C(CTRL_IDEC1_cu_system_inst_bF_buf6), .Q(_246_) );
ON21X1 ON21X1_66 ( .gnd!(gnd!), .vdd!(vdd!), .A(_245_), .B(_246_), .C(_244_), .Q(_247_) );
INX1 INX1_29 ( .gnd!(gnd!), .vdd!(vdd!), .A(PC_17_), .Q(_248_) );
ON21X1 ON21X1_67 ( .gnd!(gnd!), .vdd!(vdd!), .A(_23__bF_buf2), .B(_248_), .C(_29__bF_buf6), .Q(_249_) );
AN21X1 AN21X1_25 ( .gnd!(gnd!), .vdd!(vdd!), .A(_247_), .B(_23__bF_buf5), .C(_249_), .Q(_250_) );
ON21X1 ON21X1_68 ( .gnd!(gnd!), .vdd!(vdd!), .A(_29__bF_buf3), .B(I1_17_), .C(_32__bF_buf4), .Q(_251_) );
ON21X1 ON21X1_69 ( .gnd!(gnd!), .vdd!(vdd!), .A(_250_), .B(_251_), .C(_243_), .Q(_252_) );
NA2X1 NA2X1_70 ( .gnd!(gnd!), .vdd!(vdd!), .A(_252_), .B(CTRL_cu_r2_src_bF_buf1), .Q(_253_) );
AN31X1 AN31X1_11 ( .gnd!(gnd!), .vdd!(vdd!), .A(_36__bF_buf2), .B(rfRS2[17]), .C(_39__bF_buf4), .D(_21__bF_buf0), .Q(_254_) );
AN22X1 AN22X1_11 ( .gnd!(gnd!), .vdd!(vdd!), .A(_21__bF_buf0), .B(_242_), .C(_253_), .D(_254_), .Q(_4__17_) );
INX1 INX1_30 ( .gnd!(gnd!), .vdd!(vdd!), .A(_678__18_), .Q(_255_) );
NA2X1 NA2X1_71 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_IDEC1_cu_load_inst_bF_buf3), .B(EXT_do_18_), .Q(_256_) );
NA2I1X1 NA2I1X1_19 ( .gnd!(gnd!), .vdd!(vdd!), .AN(CTRL_IDEC1_cu_system_inst_bF_buf3), .B(R_18_), .Q(_257_) );
NO2I1X1 NO2I1X1_19 ( .gnd!(gnd!), .vdd!(vdd!), .AN(CTRL_cu_csr_rd_s1_bF_buf7), .B(CNTR_Timer_18_), .Q(_258_) );
ON21X1 ON21X1_70 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_cu_csr_rd_s1_bF_buf6), .B(CNTR_Cycle_18_), .C(CTRL_IDEC1_cu_system_inst_bF_buf2), .Q(_259_) );
ON21X1 ON21X1_71 ( .gnd!(gnd!), .vdd!(vdd!), .A(_258_), .B(_259_), .C(_257_), .Q(_260_) );
INX1 INX1_31 ( .gnd!(gnd!), .vdd!(vdd!), .A(PC_18_), .Q(_261_) );
ON21X1 ON21X1_72 ( .gnd!(gnd!), .vdd!(vdd!), .A(_23__bF_buf2), .B(_261_), .C(_29__bF_buf6), .Q(_262_) );
AN21X1 AN21X1_26 ( .gnd!(gnd!), .vdd!(vdd!), .A(_260_), .B(_23__bF_buf2), .C(_262_), .Q(_263_) );
ON21X1 ON21X1_73 ( .gnd!(gnd!), .vdd!(vdd!), .A(_29__bF_buf4), .B(I1_18_), .C(_32__bF_buf0), .Q(_264_) );
ON21X1 ON21X1_74 ( .gnd!(gnd!), .vdd!(vdd!), .A(_263_), .B(_264_), .C(_256_), .Q(_265_) );
NA2X1 NA2X1_72 ( .gnd!(gnd!), .vdd!(vdd!), .A(_265_), .B(CTRL_cu_r2_src_bF_buf3), .Q(_266_) );
AN31X1 AN31X1_12 ( .gnd!(gnd!), .vdd!(vdd!), .A(_36__bF_buf0), .B(rfRS2[18]), .C(_39__bF_buf2), .D(_21__bF_buf1), .Q(_267_) );
AN22X1 AN22X1_12 ( .gnd!(gnd!), .vdd!(vdd!), .A(_21__bF_buf1), .B(_255_), .C(_266_), .D(_267_), .Q(_4__18_) );
INX1 INX1_32 ( .gnd!(gnd!), .vdd!(vdd!), .A(_678__19_), .Q(_269_) );
NA2X1 NA2X1_73 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_IDEC1_cu_load_inst_bF_buf4), .B(EXT_do_19_), .Q(_270_) );
NA2I1X1 NA2I1X1_20 ( .gnd!(gnd!), .vdd!(vdd!), .AN(CTRL_IDEC1_cu_system_inst_bF_buf7), .B(R_19_), .Q(_271_) );
NO2I1X1 NO2I1X1_20 ( .gnd!(gnd!), .vdd!(vdd!), .AN(CTRL_cu_csr_rd_s1_bF_buf1), .B(CNTR_Timer_19_), .Q(_272_) );
ON21X1 ON21X1_75 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_cu_csr_rd_s1_bF_buf1), .B(CNTR_Cycle_19_), .C(CTRL_IDEC1_cu_system_inst_bF_buf5), .Q(_273_) );
ON21X1 ON21X1_76 ( .gnd!(gnd!), .vdd!(vdd!), .A(_272_), .B(_273_), .C(_271_), .Q(_274_) );
INX1 INX1_33 ( .gnd!(gnd!), .vdd!(vdd!), .A(PC_19_), .Q(_275_) );
ON21X1 ON21X1_77 ( .gnd!(gnd!), .vdd!(vdd!), .A(_23__bF_buf5), .B(_275_), .C(_29__bF_buf6), .Q(_276_) );
AN21X1 AN21X1_27 ( .gnd!(gnd!), .vdd!(vdd!), .A(_274_), .B(_23__bF_buf4), .C(_276_), .Q(_277_) );
ON21X1 ON21X1_78 ( .gnd!(gnd!), .vdd!(vdd!), .A(_29__bF_buf2), .B(I1_19_), .C(_32__bF_buf0), .Q(_278_) );
ON21X1 ON21X1_79 ( .gnd!(gnd!), .vdd!(vdd!), .A(_277_), .B(_278_), .C(_270_), .Q(_279_) );
NA2X1 NA2X1_74 ( .gnd!(gnd!), .vdd!(vdd!), .A(_279_), .B(CTRL_cu_r2_src_bF_buf4), .Q(_280_) );
AN31X1 AN31X1_13 ( .gnd!(gnd!), .vdd!(vdd!), .A(_36__bF_buf3), .B(rfRS2[19]), .C(_39__bF_buf1), .D(_21__bF_buf7), .Q(_281_) );
AN22X1 AN22X1_13 ( .gnd!(gnd!), .vdd!(vdd!), .A(_21__bF_buf2), .B(_269_), .C(_280_), .D(_281_), .Q(_4__19_) );
NA2X1 NA2X1_75 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_IDEC1_cu_load_inst_bF_buf1), .B(EXT_do_20_), .Q(_282_) );
NA2I1X1 NA2I1X1_21 ( .gnd!(gnd!), .vdd!(vdd!), .AN(CTRL_IDEC1_cu_system_inst_bF_buf7), .B(R_20_), .Q(_283_) );
NO2I1X1 NO2I1X1_21 ( .gnd!(gnd!), .vdd!(vdd!), .AN(CTRL_cu_csr_rd_s1_bF_buf7), .B(CNTR_Timer_20_), .Q(_284_) );
ON21X1 ON21X1_80 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_cu_csr_rd_s1_bF_buf7), .B(CNTR_Cycle_20_), .C(CTRL_IDEC1_cu_system_inst_bF_buf2), .Q(_285_) );
ON211X1 ON211X1_15 ( .gnd!(gnd!), .vdd!(vdd!), .A(_284_), .B(_285_), .C(_23__bF_buf4), .D(_283_), .Q(_286_) );
INX1 INX1_34 ( .gnd!(gnd!), .vdd!(vdd!), .A(PC_20_), .Q(_287_) );
NA2X1 NA2X1_76 ( .gnd!(gnd!), .vdd!(vdd!), .A(_287_), .B(CTRL_cu_j_inst_1), .Q(_288_) );
AN21X1 AN21X1_28 ( .gnd!(gnd!), .vdd!(vdd!), .A(_286_), .B(_288_), .C(CTRL_IDEC1_cu_lui_inst), .Q(_289_) );
ON21X1 ON21X1_81 ( .gnd!(gnd!), .vdd!(vdd!), .A(_29__bF_buf3), .B(I1_20_), .C(_32__bF_buf4), .Q(_290_) );
ON211X1 ON211X1_16 ( .gnd!(gnd!), .vdd!(vdd!), .A(_289_), .B(_290_), .C(CTRL_cu_r2_src_bF_buf5), .D(_282_), .Q(_291_) );
AN21X1 AN21X1_29 ( .gnd!(gnd!), .vdd!(vdd!), .A(_39__bF_buf1), .B(rfRS2[20]), .C(CTRL_cu_r2_src_bF_buf0), .Q(_292_) );
NO2X1 NO2X1_72 ( .gnd!(gnd!), .vdd!(vdd!), .A(_21__bF_buf6), .B(_292_), .Q(_293_) );
AO22X2 AO22X2_8 ( .gnd!(gnd!), .vdd!(vdd!), .A(_21__bF_buf6), .B(_678__20_), .C(_291_), .D(_293_), .Q(_4__20_) );
NA2X1 NA2X1_77 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_IDEC1_cu_load_inst_bF_buf2), .B(EXT_do_21_), .Q(_294_) );
NA2I1X1 NA2I1X1_22 ( .gnd!(gnd!), .vdd!(vdd!), .AN(CTRL_IDEC1_cu_system_inst_bF_buf6), .B(R_21_), .Q(_295_) );
NO2I1X1 NO2I1X1_22 ( .gnd!(gnd!), .vdd!(vdd!), .AN(CTRL_cu_csr_rd_s1_bF_buf4), .B(CNTR_Timer_21_), .Q(_296_) );
ON21X1 ON21X1_82 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_cu_csr_rd_s1_bF_buf7), .B(CNTR_Cycle_21_), .C(CTRL_IDEC1_cu_system_inst_bF_buf2), .Q(_297_) );
ON211X1 ON211X1_17 ( .gnd!(gnd!), .vdd!(vdd!), .A(_296_), .B(_297_), .C(_23__bF_buf4), .D(_295_), .Q(_298_) );
INX1 INX1_35 ( .gnd!(gnd!), .vdd!(vdd!), .A(PC_21_), .Q(_299_) );
NA2X1 NA2X1_78 ( .gnd!(gnd!), .vdd!(vdd!), .A(_299_), .B(CTRL_cu_j_inst_1), .Q(_300_) );
AN21X1 AN21X1_30 ( .gnd!(gnd!), .vdd!(vdd!), .A(_298_), .B(_300_), .C(CTRL_IDEC1_cu_lui_inst), .Q(_301_) );
ON21X1 ON21X1_83 ( .gnd!(gnd!), .vdd!(vdd!), .A(_29__bF_buf0), .B(I1_21_), .C(_32__bF_buf3), .Q(_302_) );
ON211X1 ON211X1_18 ( .gnd!(gnd!), .vdd!(vdd!), .A(_301_), .B(_302_), .C(CTRL_cu_r2_src_bF_buf2), .D(_294_), .Q(_303_) );
AN21X1 AN21X1_31 ( .gnd!(gnd!), .vdd!(vdd!), .A(_39__bF_buf0), .B(rfRS2[21]), .C(CTRL_cu_r2_src_bF_buf0), .Q(_304_) );
NO2X1 NO2X1_73 ( .gnd!(gnd!), .vdd!(vdd!), .A(_21__bF_buf7), .B(_304_), .Q(_305_) );
AO22X2 AO22X2_9 ( .gnd!(gnd!), .vdd!(vdd!), .A(_21__bF_buf6), .B(_678__21_), .C(_303_), .D(_305_), .Q(_4__21_) );
INX1 INX1_36 ( .gnd!(gnd!), .vdd!(vdd!), .A(_678__22_), .Q(_306_) );
NA2X1 NA2X1_79 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_IDEC1_cu_load_inst_bF_buf4), .B(EXT_do_22_), .Q(_307_) );
NA2I1X1 NA2I1X1_23 ( .gnd!(gnd!), .vdd!(vdd!), .AN(CTRL_IDEC1_cu_system_inst_bF_buf7), .B(R_22_), .Q(_308_) );
NO2I1X1 NO2I1X1_23 ( .gnd!(gnd!), .vdd!(vdd!), .AN(CTRL_cu_csr_rd_s1_bF_buf3), .B(CNTR_Timer_22_), .Q(_309_) );
ON21X1 ON21X1_84 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_cu_csr_rd_s1_bF_buf3), .B(CNTR_Cycle_22_), .C(CTRL_IDEC1_cu_system_inst_bF_buf2), .Q(_310_) );
ON21X1 ON21X1_85 ( .gnd!(gnd!), .vdd!(vdd!), .A(_309_), .B(_310_), .C(_308_), .Q(_311_) );
INX1 INX1_37 ( .gnd!(gnd!), .vdd!(vdd!), .A(PC_22_), .Q(_312_) );
ON21X1 ON21X1_86 ( .gnd!(gnd!), .vdd!(vdd!), .A(_23__bF_buf3), .B(_312_), .C(_29__bF_buf4), .Q(_313_) );
AN21X1 AN21X1_32 ( .gnd!(gnd!), .vdd!(vdd!), .A(_311_), .B(_23__bF_buf3), .C(_313_), .Q(_314_) );
ON21X1 ON21X1_87 ( .gnd!(gnd!), .vdd!(vdd!), .A(_29__bF_buf4), .B(I1_22_), .C(_32__bF_buf0), .Q(_315_) );
ON21X1 ON21X1_88 ( .gnd!(gnd!), .vdd!(vdd!), .A(_314_), .B(_315_), .C(_307_), .Q(_316_) );
NA2X1 NA2X1_80 ( .gnd!(gnd!), .vdd!(vdd!), .A(_316_), .B(CTRL_cu_r2_src_bF_buf1), .Q(_317_) );
AN31X1 AN31X1_14 ( .gnd!(gnd!), .vdd!(vdd!), .A(_36__bF_buf2), .B(rfRS2[22]), .C(_39__bF_buf4), .D(_21__bF_buf0), .Q(_318_) );
AN22X1 AN22X1_14 ( .gnd!(gnd!), .vdd!(vdd!), .A(_21__bF_buf0), .B(_306_), .C(_317_), .D(_318_), .Q(_4__22_) );
INX1 INX1_38 ( .gnd!(gnd!), .vdd!(vdd!), .A(_678__23_), .Q(_319_) );
NA2X1 NA2X1_81 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_IDEC1_cu_load_inst_bF_buf3), .B(EXT_do_23_), .Q(_320_) );
NA2I1X1 NA2I1X1_24 ( .gnd!(gnd!), .vdd!(vdd!), .AN(CTRL_IDEC1_cu_system_inst_bF_buf0), .B(R_23_), .Q(_321_) );
NO2I1X1 NO2I1X1_24 ( .gnd!(gnd!), .vdd!(vdd!), .AN(CTRL_cu_csr_rd_s1_bF_buf5), .B(CNTR_Timer_23_), .Q(_322_) );
ON21X1 ON21X1_89 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_cu_csr_rd_s1_bF_buf6), .B(CNTR_Cycle_23_), .C(CTRL_IDEC1_cu_system_inst_bF_buf1), .Q(_323_) );
ON21X1 ON21X1_90 ( .gnd!(gnd!), .vdd!(vdd!), .A(_322_), .B(_323_), .C(_321_), .Q(_324_) );
INX1 INX1_39 ( .gnd!(gnd!), .vdd!(vdd!), .A(PC_23_), .Q(_325_) );
ON21X1 ON21X1_91 ( .gnd!(gnd!), .vdd!(vdd!), .A(_23__bF_buf6), .B(_325_), .C(_29__bF_buf5), .Q(_326_) );
AN21X1 AN21X1_33 ( .gnd!(gnd!), .vdd!(vdd!), .A(_324_), .B(_23__bF_buf3), .C(_326_), .Q(_327_) );
ON21X1 ON21X1_92 ( .gnd!(gnd!), .vdd!(vdd!), .A(_29__bF_buf3), .B(I1_23_), .C(_32__bF_buf4), .Q(_328_) );
ON21X1 ON21X1_93 ( .gnd!(gnd!), .vdd!(vdd!), .A(_327_), .B(_328_), .C(_320_), .Q(_329_) );
NA2X1 NA2X1_82 ( .gnd!(gnd!), .vdd!(vdd!), .A(_329_), .B(CTRL_cu_r2_src_bF_buf0), .Q(_330_) );
AN31X1 AN31X1_15 ( .gnd!(gnd!), .vdd!(vdd!), .A(_36__bF_buf2), .B(rfRS2[23]), .C(_39__bF_buf4), .D(_21__bF_buf0), .Q(_331_) );
AN22X1 AN22X1_15 ( .gnd!(gnd!), .vdd!(vdd!), .A(_21__bF_buf0), .B(_319_), .C(_330_), .D(_331_), .Q(_4__23_) );
INX1 INX1_40 ( .gnd!(gnd!), .vdd!(vdd!), .A(_678__24_), .Q(_332_) );
NA2X1 NA2X1_83 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_IDEC1_cu_load_inst_bF_buf3), .B(EXT_do_24_), .Q(_333_) );
NA2I1X1 NA2I1X1_25 ( .gnd!(gnd!), .vdd!(vdd!), .AN(CTRL_IDEC1_cu_system_inst_bF_buf7), .B(R_24_), .Q(_334_) );
NO2I1X1 NO2I1X1_25 ( .gnd!(gnd!), .vdd!(vdd!), .AN(CTRL_cu_csr_rd_s1_bF_buf4), .B(CNTR_Timer_24_), .Q(_335_) );
ON21X1 ON21X1_94 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_cu_csr_rd_s1_bF_buf7), .B(CNTR_Cycle_24_), .C(CTRL_IDEC1_cu_system_inst_bF_buf2), .Q(_336_) );
ON21X1 ON21X1_95 ( .gnd!(gnd!), .vdd!(vdd!), .A(_335_), .B(_336_), .C(_334_), .Q(_337_) );
INX1 INX1_41 ( .gnd!(gnd!), .vdd!(vdd!), .A(PC_24_), .Q(_338_) );
ON21X1 ON21X1_96 ( .gnd!(gnd!), .vdd!(vdd!), .A(_23__bF_buf1), .B(_338_), .C(_29__bF_buf2), .Q(_339_) );
AN21X1 AN21X1_34 ( .gnd!(gnd!), .vdd!(vdd!), .A(_337_), .B(_23__bF_buf1), .C(_339_), .Q(_340_) );
ON21X1 ON21X1_97 ( .gnd!(gnd!), .vdd!(vdd!), .A(_29__bF_buf5), .B(I1_24_), .C(_32__bF_buf2), .Q(_341_) );
ON21X1 ON21X1_98 ( .gnd!(gnd!), .vdd!(vdd!), .A(_340_), .B(_341_), .C(_333_), .Q(_342_) );
NA2X1 NA2X1_84 ( .gnd!(gnd!), .vdd!(vdd!), .A(_342_), .B(CTRL_cu_r2_src_bF_buf2), .Q(_343_) );
AN31X1 AN31X1_16 ( .gnd!(gnd!), .vdd!(vdd!), .A(_36__bF_buf3), .B(rfRS2[24]), .C(_39__bF_buf1), .D(_21__bF_buf3), .Q(_344_) );
AN22X1 AN22X1_16 ( .gnd!(gnd!), .vdd!(vdd!), .A(_21__bF_buf3), .B(_332_), .C(_343_), .D(_344_), .Q(_4__24_) );
INX1 INX1_42 ( .gnd!(gnd!), .vdd!(vdd!), .A(_678__25_), .Q(_345_) );
NA2X1 NA2X1_85 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_IDEC1_cu_load_inst_bF_buf0), .B(EXT_do_25_), .Q(_346_) );
NA2I1X1 NA2I1X1_26 ( .gnd!(gnd!), .vdd!(vdd!), .AN(CTRL_IDEC1_cu_system_inst_bF_buf3), .B(R_25_), .Q(_347_) );
NO2I1X1 NO2I1X1_26 ( .gnd!(gnd!), .vdd!(vdd!), .AN(CTRL_cu_csr_rd_s1_bF_buf4), .B(CNTR_Timer_25_), .Q(_348_) );
ON21X1 ON21X1_99 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_cu_csr_rd_s1_bF_buf7), .B(CNTR_Cycle_25_), .C(CTRL_IDEC1_cu_system_inst_bF_buf6), .Q(_349_) );
ON21X1 ON21X1_100 ( .gnd!(gnd!), .vdd!(vdd!), .A(_348_), .B(_349_), .C(_347_), .Q(_350_) );
INX1 INX1_43 ( .gnd!(gnd!), .vdd!(vdd!), .A(PC_25_), .Q(_351_) );
ON21X1 ON21X1_101 ( .gnd!(gnd!), .vdd!(vdd!), .A(_23__bF_buf6), .B(_351_), .C(_29__bF_buf5), .Q(_352_) );
AN21X1 AN21X1_35 ( .gnd!(gnd!), .vdd!(vdd!), .A(_350_), .B(_23__bF_buf6), .C(_352_), .Q(_353_) );
ON21X1 ON21X1_102 ( .gnd!(gnd!), .vdd!(vdd!), .A(_29__bF_buf3), .B(I1_25_), .C(_32__bF_buf4), .Q(_354_) );
ON21X1 ON21X1_103 ( .gnd!(gnd!), .vdd!(vdd!), .A(_353_), .B(_354_), .C(_346_), .Q(_355_) );
NA2X1 NA2X1_86 ( .gnd!(gnd!), .vdd!(vdd!), .A(_355_), .B(CTRL_cu_r2_src_bF_buf2), .Q(_356_) );
AN31X1 AN31X1_17 ( .gnd!(gnd!), .vdd!(vdd!), .A(_36__bF_buf3), .B(rfRS2[25]), .C(_39__bF_buf1), .D(_21__bF_buf3), .Q(_357_) );
AN22X1 AN22X1_17 ( .gnd!(gnd!), .vdd!(vdd!), .A(_21__bF_buf3), .B(_345_), .C(_356_), .D(_357_), .Q(_4__25_) );
INX1 INX1_44 ( .gnd!(gnd!), .vdd!(vdd!), .A(_678__26_), .Q(_358_) );
NA2X1 NA2X1_87 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_IDEC1_cu_load_inst_bF_buf2), .B(EXT_do_26_), .Q(_359_) );
NA2I1X1 NA2I1X1_27 ( .gnd!(gnd!), .vdd!(vdd!), .AN(CTRL_IDEC1_cu_system_inst_bF_buf0), .B(R_26_), .Q(_360_) );
NO2I1X1 NO2I1X1_27 ( .gnd!(gnd!), .vdd!(vdd!), .AN(CTRL_cu_csr_rd_s1_bF_buf4), .B(CNTR_Timer_26_), .Q(_361_) );
ON21X1 ON21X1_104 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_cu_csr_rd_s1_bF_buf6), .B(CNTR_Cycle_26_), .C(CTRL_IDEC1_cu_system_inst_bF_buf1), .Q(_362_) );
ON21X1 ON21X1_105 ( .gnd!(gnd!), .vdd!(vdd!), .A(_361_), .B(_362_), .C(_360_), .Q(_363_) );
INX1 INX1_45 ( .gnd!(gnd!), .vdd!(vdd!), .A(PC_26_), .Q(_364_) );
ON21X1 ON21X1_106 ( .gnd!(gnd!), .vdd!(vdd!), .A(_23__bF_buf3), .B(_364_), .C(_29__bF_buf4), .Q(_365_) );
AN21X1 AN21X1_36 ( .gnd!(gnd!), .vdd!(vdd!), .A(_363_), .B(_23__bF_buf6), .C(_365_), .Q(_366_) );
ON21X1 ON21X1_107 ( .gnd!(gnd!), .vdd!(vdd!), .A(_29__bF_buf3), .B(I1_26_), .C(_32__bF_buf4), .Q(_367_) );
ON21X1 ON21X1_108 ( .gnd!(gnd!), .vdd!(vdd!), .A(_366_), .B(_367_), .C(_359_), .Q(_368_) );
NA2X1 NA2X1_88 ( .gnd!(gnd!), .vdd!(vdd!), .A(_368_), .B(CTRL_cu_r2_src_bF_buf0), .Q(_369_) );
AN31X1 AN31X1_18 ( .gnd!(gnd!), .vdd!(vdd!), .A(_36__bF_buf0), .B(rfRS2[26]), .C(_39__bF_buf2), .D(_21__bF_buf7), .Q(_370_) );
AN22X1 AN22X1_18 ( .gnd!(gnd!), .vdd!(vdd!), .A(_21__bF_buf7), .B(_358_), .C(_369_), .D(_370_), .Q(_4__26_) );
NA2X1 NA2X1_89 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_IDEC1_cu_load_inst_bF_buf4), .B(EXT_do_27_), .Q(_371_) );
NA2I1X1 NA2I1X1_28 ( .gnd!(gnd!), .vdd!(vdd!), .AN(CTRL_IDEC1_cu_system_inst_bF_buf0), .B(R_27_), .Q(_372_) );
NO2I1X1 NO2I1X1_28 ( .gnd!(gnd!), .vdd!(vdd!), .AN(CTRL_cu_csr_rd_s1_bF_buf3), .B(CNTR_Timer_27_), .Q(_373_) );
ON21X1 ON21X1_109 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_cu_csr_rd_s1_bF_buf6), .B(CNTR_Cycle_27_), .C(CTRL_IDEC1_cu_system_inst_bF_buf1), .Q(_374_) );
ON211X1 ON211X1_19 ( .gnd!(gnd!), .vdd!(vdd!), .A(_373_), .B(_374_), .C(_23__bF_buf0), .D(_372_), .Q(_375_) );
INX1 INX1_46 ( .gnd!(gnd!), .vdd!(vdd!), .A(PC_27_), .Q(_376_) );
NA2X1 NA2X1_90 ( .gnd!(gnd!), .vdd!(vdd!), .A(_376_), .B(CTRL_cu_j_inst_1), .Q(_377_) );
AN21X1 AN21X1_37 ( .gnd!(gnd!), .vdd!(vdd!), .A(_375_), .B(_377_), .C(CTRL_IDEC1_cu_lui_inst), .Q(_378_) );
ON21X1 ON21X1_110 ( .gnd!(gnd!), .vdd!(vdd!), .A(_29__bF_buf5), .B(I1_27_), .C(_32__bF_buf2), .Q(_379_) );
ON211X1 ON211X1_20 ( .gnd!(gnd!), .vdd!(vdd!), .A(_378_), .B(_379_), .C(CTRL_cu_r2_src_bF_buf5), .D(_371_), .Q(_380_) );
AN21X1 AN21X1_38 ( .gnd!(gnd!), .vdd!(vdd!), .A(_39__bF_buf2), .B(rfRS2[27]), .C(CTRL_cu_r2_src_bF_buf1), .Q(_381_) );
NO2X1 NO2X1_74 ( .gnd!(gnd!), .vdd!(vdd!), .A(_21__bF_buf7), .B(_381_), .Q(_382_) );
AO22X2 AO22X2_10 ( .gnd!(gnd!), .vdd!(vdd!), .A(_21__bF_buf7), .B(_678__27_), .C(_380_), .D(_382_), .Q(_4__27_) );
NA2X1 NA2X1_91 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_IDEC1_cu_load_inst_bF_buf1), .B(EXT_do_28_), .Q(_383_) );
NA2I1X1 NA2I1X1_29 ( .gnd!(gnd!), .vdd!(vdd!), .AN(CTRL_IDEC1_cu_system_inst_bF_buf6), .B(R_28_), .Q(_384_) );
NO2I1X1 NO2I1X1_29 ( .gnd!(gnd!), .vdd!(vdd!), .AN(CTRL_cu_csr_rd_s1_bF_buf4), .B(CNTR_Timer_28_), .Q(_385_) );
ON21X1 ON21X1_111 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_cu_csr_rd_s1_bF_buf6), .B(CNTR_Cycle_28_), .C(CTRL_IDEC1_cu_system_inst_bF_buf1), .Q(_386_) );
ON211X1 ON211X1_21 ( .gnd!(gnd!), .vdd!(vdd!), .A(_385_), .B(_386_), .C(_23__bF_buf0), .D(_384_), .Q(_387_) );
INX1 INX1_47 ( .gnd!(gnd!), .vdd!(vdd!), .A(PC_28_), .Q(_388_) );
NA2X1 NA2X1_92 ( .gnd!(gnd!), .vdd!(vdd!), .A(_388_), .B(CTRL_cu_j_inst_1), .Q(_389_) );
AN21X1 AN21X1_39 ( .gnd!(gnd!), .vdd!(vdd!), .A(_387_), .B(_389_), .C(CTRL_IDEC1_cu_lui_inst), .Q(_390_) );
ON21X1 ON21X1_112 ( .gnd!(gnd!), .vdd!(vdd!), .A(_29__bF_buf0), .B(I1_28_), .C(_32__bF_buf3), .Q(_391_) );
ON211X1 ON211X1_22 ( .gnd!(gnd!), .vdd!(vdd!), .A(_390_), .B(_391_), .C(CTRL_cu_r2_src_bF_buf5), .D(_383_), .Q(_392_) );
AN21X1 AN21X1_40 ( .gnd!(gnd!), .vdd!(vdd!), .A(_39__bF_buf0), .B(rfRS2[28]), .C(CTRL_cu_r2_src_bF_buf0), .Q(_393_) );
NO2X1 NO2X1_75 ( .gnd!(gnd!), .vdd!(vdd!), .A(_21__bF_buf6), .B(_393_), .Q(_394_) );
AO22X2 AO22X2_11 ( .gnd!(gnd!), .vdd!(vdd!), .A(_21__bF_buf6), .B(_678__28_), .C(_392_), .D(_394_), .Q(_4__28_) );
INX1 INX1_48 ( .gnd!(gnd!), .vdd!(vdd!), .A(_678__29_), .Q(_395_) );
NA2X1 NA2X1_93 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_IDEC1_cu_load_inst_bF_buf3), .B(EXT_do_29_), .Q(_396_) );
NA2I1X1 NA2I1X1_30 ( .gnd!(gnd!), .vdd!(vdd!), .AN(CTRL_IDEC1_cu_system_inst_bF_buf7), .B(R_29_), .Q(_397_) );
NO2I1X1 NO2I1X1_30 ( .gnd!(gnd!), .vdd!(vdd!), .AN(CTRL_cu_csr_rd_s1_bF_buf4), .B(CNTR_Timer_29_), .Q(_398_) );
ON21X1 ON21X1_113 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_cu_csr_rd_s1_bF_buf6), .B(CNTR_Cycle_29_), .C(CTRL_IDEC1_cu_system_inst_bF_buf2), .Q(_399_) );
ON21X1 ON21X1_114 ( .gnd!(gnd!), .vdd!(vdd!), .A(_398_), .B(_399_), .C(_397_), .Q(_400_) );
INX1 INX1_49 ( .gnd!(gnd!), .vdd!(vdd!), .A(PC_29_), .Q(_401_) );
ON21X1 ON21X1_115 ( .gnd!(gnd!), .vdd!(vdd!), .A(_23__bF_buf2), .B(_401_), .C(_29__bF_buf6), .Q(_402_) );
AN21X1 AN21X1_41 ( .gnd!(gnd!), .vdd!(vdd!), .A(_400_), .B(_23__bF_buf2), .C(_402_), .Q(_403_) );
ON21X1 ON21X1_116 ( .gnd!(gnd!), .vdd!(vdd!), .A(_29__bF_buf3), .B(I1_29_), .C(_32__bF_buf4), .Q(_404_) );
ON21X1 ON21X1_117 ( .gnd!(gnd!), .vdd!(vdd!), .A(_403_), .B(_404_), .C(_396_), .Q(_405_) );
NA2X1 NA2X1_94 ( .gnd!(gnd!), .vdd!(vdd!), .A(_405_), .B(CTRL_cu_r2_src_bF_buf4), .Q(_406_) );
AN31X1 AN31X1_19 ( .gnd!(gnd!), .vdd!(vdd!), .A(_36__bF_buf1), .B(rfRS2[29]), .C(_39__bF_buf2), .D(_21__bF_buf1), .Q(_407_) );
AN22X1 AN22X1_19 ( .gnd!(gnd!), .vdd!(vdd!), .A(_21__bF_buf2), .B(_395_), .C(_406_), .D(_407_), .Q(_4__29_) );
INX1 INX1_50 ( .gnd!(gnd!), .vdd!(vdd!), .A(_678__30_), .Q(_408_) );
NA2X1 NA2X1_95 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_IDEC1_cu_load_inst_bF_buf0), .B(EXT_do_30_), .Q(_409_) );
NA2I1X1 NA2I1X1_31 ( .gnd!(gnd!), .vdd!(vdd!), .AN(CTRL_IDEC1_cu_system_inst_bF_buf0), .B(R_30_), .Q(_410_) );
NO2I1X1 NO2I1X1_31 ( .gnd!(gnd!), .vdd!(vdd!), .AN(CTRL_cu_csr_rd_s1_bF_buf5), .B(CNTR_Timer_30_), .Q(_411_) );
ON21X1 ON21X1_118 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_cu_csr_rd_s1_bF_buf6), .B(CNTR_Cycle_30_), .C(CTRL_IDEC1_cu_system_inst_bF_buf1), .Q(_412_) );
ON21X1 ON21X1_119 ( .gnd!(gnd!), .vdd!(vdd!), .A(_411_), .B(_412_), .C(_410_), .Q(_413_) );
INX1 INX1_51 ( .gnd!(gnd!), .vdd!(vdd!), .A(PC_30_), .Q(_414_) );
ON21X1 ON21X1_120 ( .gnd!(gnd!), .vdd!(vdd!), .A(_23__bF_buf6), .B(_414_), .C(_29__bF_buf3), .Q(_415_) );
AN21X1 AN21X1_42 ( .gnd!(gnd!), .vdd!(vdd!), .A(_413_), .B(_23__bF_buf6), .C(_415_), .Q(_416_) );
ON21X1 ON21X1_121 ( .gnd!(gnd!), .vdd!(vdd!), .A(_29__bF_buf3), .B(I1_30_), .C(_32__bF_buf4), .Q(_417_) );
ON21X1 ON21X1_122 ( .gnd!(gnd!), .vdd!(vdd!), .A(_416_), .B(_417_), .C(_409_), .Q(_418_) );
NA2X1 NA2X1_96 ( .gnd!(gnd!), .vdd!(vdd!), .A(_418_), .B(CTRL_cu_r2_src_bF_buf4), .Q(_419_) );
AN31X1 AN31X1_20 ( .gnd!(gnd!), .vdd!(vdd!), .A(_36__bF_buf3), .B(rfRS2[30]), .C(_39__bF_buf1), .D(_21__bF_buf3), .Q(_420_) );
AN22X1 AN22X1_20 ( .gnd!(gnd!), .vdd!(vdd!), .A(_21__bF_buf7), .B(_408_), .C(_419_), .D(_420_), .Q(_4__30_) );
INX1 INX1_52 ( .gnd!(gnd!), .vdd!(vdd!), .A(_678__31_), .Q(_421_) );
NA2X1 NA2X1_97 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_IDEC1_cu_load_inst_bF_buf4), .B(EXT_do_31_), .Q(_422_) );
NA2I1X1 NA2I1X1_32 ( .gnd!(gnd!), .vdd!(vdd!), .AN(CTRL_IDEC1_cu_system_inst_bF_buf3), .B(R_31_), .Q(_423_) );
NO2I1X1 NO2I1X1_32 ( .gnd!(gnd!), .vdd!(vdd!), .AN(CTRL_cu_csr_rd_s1_bF_buf1), .B(CNTR_Timer_31_), .Q(_424_) );
ON21X1 ON21X1_123 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_cu_csr_rd_s1_bF_buf1), .B(CNTR_Cycle_31_), .C(CTRL_IDEC1_cu_system_inst_bF_buf5), .Q(_425_) );
ON21X1 ON21X1_124 ( .gnd!(gnd!), .vdd!(vdd!), .A(_424_), .B(_425_), .C(_423_), .Q(_426_) );
INX1 INX1_53 ( .gnd!(gnd!), .vdd!(vdd!), .A(PC_31_), .Q(_427_) );
ON21X1 ON21X1_125 ( .gnd!(gnd!), .vdd!(vdd!), .A(_23__bF_buf2), .B(_427_), .C(_29__bF_buf6), .Q(_428_) );
AN21X1 AN21X1_43 ( .gnd!(gnd!), .vdd!(vdd!), .A(_426_), .B(_23__bF_buf2), .C(_428_), .Q(_429_) );
ON21X1 ON21X1_126 ( .gnd!(gnd!), .vdd!(vdd!), .A(_29__bF_buf6), .B(I1_31_), .C(_32__bF_buf0), .Q(_430_) );
ON21X1 ON21X1_127 ( .gnd!(gnd!), .vdd!(vdd!), .A(_429_), .B(_430_), .C(_422_), .Q(_431_) );
NA2X1 NA2X1_98 ( .gnd!(gnd!), .vdd!(vdd!), .A(_431_), .B(CTRL_cu_r2_src_bF_buf4), .Q(_432_) );
AN31X1 AN31X1_21 ( .gnd!(gnd!), .vdd!(vdd!), .A(_36__bF_buf0), .B(rfRS2[31]), .C(_39__bF_buf2), .D(_21__bF_buf1), .Q(_433_) );
AN22X1 AN22X1_21 ( .gnd!(gnd!), .vdd!(vdd!), .A(_21__bF_buf6), .B(_421_), .C(_432_), .D(_433_), .Q(_4__31_) );
INX2 INX2_4 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_cyc_bF_buf10_bF_buf2), .Q(_434_) );
MU2X1 MU2X1_1 ( .gnd!(gnd!), .vdd!(vdd!), .IN0(_34_), .IN1(_684__0_), .Q(_5__0_), .S(_434__bF_buf3) );
OR2X2 OR2X2_1 ( .gnd!(gnd!), .vdd!(vdd!), .A(_48_), .B(_49_), .Q(_435_) );
NO2X1 NO2X1_76 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_cyc_bF_buf9_bF_buf0), .B(_684__1_), .Q(_436_) );
AN31X1 AN31X1_22 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_cyc_bF_buf8_bF_buf1), .B(_41_), .C(_435_), .D(_436_), .Q(_5__1_) );
MU2X1 MU2X1_2 ( .gnd!(gnd!), .vdd!(vdd!), .IN0(_63_), .IN1(_684__2_), .Q(_5__2_), .S(_434__bF_buf2) );
OR2X2 OR2X2_2 ( .gnd!(gnd!), .vdd!(vdd!), .A(_73_), .B(_74_), .Q(_437_) );
NO2X1 NO2X1_77 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_cyc_bF_buf7_bF_buf0), .B(_684__3_), .Q(_438_) );
AN31X1 AN31X1_23 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_cyc_bF_buf6_bF_buf1), .B(_66_), .C(_437_), .D(_438_), .Q(_5__3_) );
MU2X1 MU2X1_3 ( .gnd!(gnd!), .vdd!(vdd!), .IN0(_88_), .IN1(_684__4_), .Q(_5__4_), .S(_434__bF_buf2) );
OR2X2 OR2X2_3 ( .gnd!(gnd!), .vdd!(vdd!), .A(_98_), .B(_99_), .Q(_439_) );
NO2X1 NO2X1_78 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_cyc_bF_buf5_bF_buf0), .B(_684__5_), .Q(_440_) );
AN31X1 AN31X1_24 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_cyc_bF_buf4_bF_buf1), .B(_91_), .C(_439_), .D(_440_), .Q(_5__5_) );
MU2X1 MU2X1_4 ( .gnd!(gnd!), .vdd!(vdd!), .IN0(_113_), .IN1(_684__6_), .Q(_5__6_), .S(_434__bF_buf1) );
OR2X2 OR2X2_4 ( .gnd!(gnd!), .vdd!(vdd!), .A(_123_), .B(_124_), .Q(_441_) );
NO2X1 NO2X1_79 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_cyc_bF_buf3_bF_buf2), .B(_684__7_), .Q(_442_) );
AN31X1 AN31X1_25 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_cyc_bF_buf2_bF_buf1), .B(_116_), .C(_441_), .D(_442_), .Q(_5__7_) );
OR2X2 OR2X2_5 ( .gnd!(gnd!), .vdd!(vdd!), .A(_135_), .B(_136_), .Q(_443_) );
NO2X1 NO2X1_80 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_cyc_bF_buf1_bF_buf2), .B(_684__8_), .Q(_444_) );
AN31X1 AN31X1_26 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_cyc_bF_buf0_bF_buf2), .B(_128_), .C(_443_), .D(_444_), .Q(_5__8_) );
MU2X1 MU2X1_5 ( .gnd!(gnd!), .vdd!(vdd!), .IN0(_150_), .IN1(_684__9_), .Q(_5__9_), .S(_434__bF_buf3) );
MU2X1 MU2X1_6 ( .gnd!(gnd!), .vdd!(vdd!), .IN0(_163_), .IN1(_684__10_), .Q(_5__10_), .S(_434__bF_buf1) );
MU2X1 MU2X1_7 ( .gnd!(gnd!), .vdd!(vdd!), .IN0(_176_), .IN1(_684__11_), .Q(_5__11_), .S(_434__bF_buf0) );
MU2X1 MU2X1_8 ( .gnd!(gnd!), .vdd!(vdd!), .IN0(_189_), .IN1(_684__12_), .Q(_5__12_), .S(_434__bF_buf3) );
OR2X2 OR2X2_6 ( .gnd!(gnd!), .vdd!(vdd!), .A(_199_), .B(_200_), .Q(_445_) );
NO2X1 NO2X1_81 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_cyc_bF_buf14_bF_buf3), .B(_684__13_), .Q(_446_) );
AN31X1 AN31X1_27 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_cyc_bF_buf13_bF_buf0), .B(_192_), .C(_445_), .D(_446_), .Q(_5__13_) );
MU2X1 MU2X1_9 ( .gnd!(gnd!), .vdd!(vdd!), .IN0(_214_), .IN1(_684__14_), .Q(_5__14_), .S(_434__bF_buf2) );
MU2X1 MU2X1_10 ( .gnd!(gnd!), .vdd!(vdd!), .IN0(_227_), .IN1(_684__15_), .Q(_5__15_), .S(_434__bF_buf0) );
OR2X2 OR2X2_7 ( .gnd!(gnd!), .vdd!(vdd!), .A(_237_), .B(_238_), .Q(_447_) );
NO2X1 NO2X1_82 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_cyc_bF_buf12_bF_buf1), .B(_684__16_), .Q(_448_) );
AN31X1 AN31X1_28 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_cyc_bF_buf11_bF_buf0), .B(_230_), .C(_447_), .D(_448_), .Q(_5__16_) );
MU2X1 MU2X1_11 ( .gnd!(gnd!), .vdd!(vdd!), .IN0(_252_), .IN1(_684__17_), .Q(_5__17_), .S(_434__bF_buf3) );
MU2X1 MU2X1_12 ( .gnd!(gnd!), .vdd!(vdd!), .IN0(_265_), .IN1(_684__18_), .Q(_5__18_), .S(_434__bF_buf2) );
MU2X1 MU2X1_13 ( .gnd!(gnd!), .vdd!(vdd!), .IN0(_279_), .IN1(_684__19_), .Q(_5__19_), .S(_434__bF_buf3) );
OR2X2 OR2X2_8 ( .gnd!(gnd!), .vdd!(vdd!), .A(_289_), .B(_290_), .Q(_449_) );
NO2X1 NO2X1_83 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_cyc_bF_buf10_bF_buf2), .B(_684__20_), .Q(_450_) );
AN31X1 AN31X1_29 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_cyc_bF_buf9_bF_buf0), .B(_282_), .C(_449_), .D(_450_), .Q(_5__20_) );
OR2X2 OR2X2_9 ( .gnd!(gnd!), .vdd!(vdd!), .A(_301_), .B(_302_), .Q(_451_) );
NO2X1 NO2X1_84 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_cyc_bF_buf8_bF_buf1), .B(_684__21_), .Q(_452_) );
AN31X1 AN31X1_30 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_cyc_bF_buf7_bF_buf0), .B(_294_), .C(_451_), .D(_452_), .Q(_5__21_) );
MU2X1 MU2X1_14 ( .gnd!(gnd!), .vdd!(vdd!), .IN0(_316_), .IN1(_684__22_), .Q(_5__22_), .S(_434__bF_buf0) );
MU2X1 MU2X1_15 ( .gnd!(gnd!), .vdd!(vdd!), .IN0(_329_), .IN1(_684__23_), .Q(_5__23_), .S(_434__bF_buf3) );
MU2X1 MU2X1_16 ( .gnd!(gnd!), .vdd!(vdd!), .IN0(_342_), .IN1(_684__24_), .Q(_5__24_), .S(_434__bF_buf1) );
MU2X1 MU2X1_17 ( .gnd!(gnd!), .vdd!(vdd!), .IN0(_355_), .IN1(_684__25_), .Q(_5__25_), .S(_434__bF_buf1) );
MU2X1 MU2X1_18 ( .gnd!(gnd!), .vdd!(vdd!), .IN0(_368_), .IN1(_684__26_), .Q(_5__26_), .S(_434__bF_buf1) );
OR2X2 OR2X2_10 ( .gnd!(gnd!), .vdd!(vdd!), .A(_378_), .B(_379_), .Q(_453_) );
NO2X1 NO2X1_85 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_cyc_bF_buf6_bF_buf0), .B(_684__27_), .Q(_454_) );
AN31X1 AN31X1_31 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_cyc_bF_buf5_bF_buf2), .B(_371_), .C(_453_), .D(_454_), .Q(_5__27_) );
OR2X2 OR2X2_11 ( .gnd!(gnd!), .vdd!(vdd!), .A(_390_), .B(_391_), .Q(_455_) );
NO2X1 NO2X1_86 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_cyc_bF_buf4_bF_buf1), .B(_684__28_), .Q(_456_) );
AN31X1 AN31X1_32 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_cyc_bF_buf3_bF_buf1), .B(_383_), .C(_455_), .D(_456_), .Q(_5__28_) );
MU2X1 MU2X1_19 ( .gnd!(gnd!), .vdd!(vdd!), .IN0(_405_), .IN1(_684__29_), .Q(_5__29_), .S(_434__bF_buf2) );
MU2X1 MU2X1_20 ( .gnd!(gnd!), .vdd!(vdd!), .IN0(_418_), .IN1(_684__30_), .Q(_5__30_), .S(_434__bF_buf0) );
MU2X1 MU2X1_21 ( .gnd!(gnd!), .vdd!(vdd!), .IN0(_431_), .IN1(_684__31_), .Q(_5__31_), .S(_434__bF_buf0) );
INX1 INX1_54 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_TMRIF), .Q(_457_) );
AN21X1 AN21X1_44 ( .gnd!(gnd!), .vdd!(vdd!), .A(_457_), .B(CTRL_cu_int_ebreak), .C(IRQ), .Q(PCU_int_vec_4_) );
NO2X1 NO2X1_87 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_TMRIF), .B(CTRL_cu_int_ebreak), .Q(_458_) );
NO2X1 NO2X1_88 ( .gnd!(gnd!), .vdd!(vdd!), .A(IRQ), .B(_458_), .Q(PCU_int_vec_5_) );
MU2X1 MU2X1_22 ( .gnd!(gnd!), .vdd!(vdd!), .IN0(_681__0_), .IN1(PC1_0_), .Q(ALU_a_0_), .S(CTRL_IDEC1_cu_auipc_inst_bF_buf2) );
MU2X1 MU2X1_23 ( .gnd!(gnd!), .vdd!(vdd!), .IN0(_681__1_), .IN1(PC1_1_), .Q(ALU_a_1_), .S(CTRL_IDEC1_cu_auipc_inst_bF_buf2) );
MU2X1 MU2X1_24 ( .gnd!(gnd!), .vdd!(vdd!), .IN0(_681__2_), .IN1(PC1_2_), .Q(ALU_a_2_), .S(CTRL_IDEC1_cu_auipc_inst_bF_buf2) );
MU2X1 MU2X1_25 ( .gnd!(gnd!), .vdd!(vdd!), .IN0(_681__3_), .IN1(PC1_3_), .Q(ALU_a_3_), .S(CTRL_IDEC1_cu_auipc_inst_bF_buf4) );
MU2X1 MU2X1_26 ( .gnd!(gnd!), .vdd!(vdd!), .IN0(_681__4_), .IN1(PC1_4_), .Q(ALU_a_4_), .S(CTRL_IDEC1_cu_auipc_inst_bF_buf1) );
INX1 INX1_55 ( .gnd!(gnd!), .vdd!(vdd!), .A(_681__5_), .Q(_459_) );
INX1 INX1_56 ( .gnd!(gnd!), .vdd!(vdd!), .A(PC1_5_), .Q(_460_) );
MU2IX1 MU2IX1_1 ( .gnd!(gnd!), .vdd!(vdd!), .IN0(_459_), .IN1(_460_), .Q(ALU_a_5_), .S(CTRL_IDEC1_cu_auipc_inst_bF_buf4) );
MU2X1 MU2X1_27 ( .gnd!(gnd!), .vdd!(vdd!), .IN0(_681__6_), .IN1(PC1_6_), .Q(ALU_a_6_), .S(CTRL_IDEC1_cu_auipc_inst_bF_buf1) );
MU2X1 MU2X1_28 ( .gnd!(gnd!), .vdd!(vdd!), .IN0(_681__7_), .IN1(PC1_7_), .Q(ALU_a_7_), .S(CTRL_IDEC1_cu_auipc_inst_bF_buf0) );
INX1 INX1_57 ( .gnd!(gnd!), .vdd!(vdd!), .A(_681__8_), .Q(_461_) );
INX1 INX1_58 ( .gnd!(gnd!), .vdd!(vdd!), .A(PC1_8_), .Q(_462_) );
MU2IX1 MU2IX1_2 ( .gnd!(gnd!), .vdd!(vdd!), .IN0(_461_), .IN1(_462_), .Q(ALU_a_8_), .S(CTRL_IDEC1_cu_auipc_inst_bF_buf1) );
MU2X1 MU2X1_29 ( .gnd!(gnd!), .vdd!(vdd!), .IN0(_681__9_), .IN1(PC1_9_), .Q(ALU_a_9_), .S(CTRL_IDEC1_cu_auipc_inst_bF_buf1) );
MU2X1 MU2X1_30 ( .gnd!(gnd!), .vdd!(vdd!), .IN0(_681__10_), .IN1(PC1_10_), .Q(ALU_a_10_), .S(CTRL_IDEC1_cu_auipc_inst_bF_buf0) );
MU2X1 MU2X1_31 ( .gnd!(gnd!), .vdd!(vdd!), .IN0(_681__11_), .IN1(PC1_11_), .Q(ALU_a_11_), .S(CTRL_IDEC1_cu_auipc_inst_bF_buf0) );
MU2X1 MU2X1_32 ( .gnd!(gnd!), .vdd!(vdd!), .IN0(_681__12_), .IN1(PC1_12_), .Q(ALU_a_12_), .S(CTRL_IDEC1_cu_auipc_inst_bF_buf0) );
MU2X1 MU2X1_33 ( .gnd!(gnd!), .vdd!(vdd!), .IN0(_681__13_), .IN1(PC1_13_), .Q(ALU_a_13_), .S(CTRL_IDEC1_cu_auipc_inst_bF_buf0) );
MU2X1 MU2X1_34 ( .gnd!(gnd!), .vdd!(vdd!), .IN0(_681__14_), .IN1(PC1_14_), .Q(ALU_a_14_), .S(CTRL_IDEC1_cu_auipc_inst_bF_buf0) );
MU2X1 MU2X1_35 ( .gnd!(gnd!), .vdd!(vdd!), .IN0(_681__15_), .IN1(PC1_15_), .Q(ALU_a_15_), .S(CTRL_IDEC1_cu_auipc_inst_bF_buf1) );
INX1 INX1_59 ( .gnd!(gnd!), .vdd!(vdd!), .A(_681__16_), .Q(_463_) );
INX1 INX1_60 ( .gnd!(gnd!), .vdd!(vdd!), .A(PC1_16_), .Q(_464_) );
MU2IX1 MU2IX1_3 ( .gnd!(gnd!), .vdd!(vdd!), .IN0(_463_), .IN1(_464_), .Q(ALU_a_16_), .S(CTRL_IDEC1_cu_auipc_inst_bF_buf1) );
MU2X1 MU2X1_36 ( .gnd!(gnd!), .vdd!(vdd!), .IN0(_681__17_), .IN1(PC1_17_), .Q(ALU_a_17_), .S(CTRL_IDEC1_cu_auipc_inst_bF_buf4) );
MU2X1 MU2X1_37 ( .gnd!(gnd!), .vdd!(vdd!), .IN0(_681__18_), .IN1(PC1_18_), .Q(ALU_a_18_), .S(CTRL_IDEC1_cu_auipc_inst_bF_buf2) );
MU2X1 MU2X1_38 ( .gnd!(gnd!), .vdd!(vdd!), .IN0(_681__19_), .IN1(PC1_19_), .Q(ALU_a_19_), .S(CTRL_IDEC1_cu_auipc_inst_bF_buf4) );
INX1 INX1_61 ( .gnd!(gnd!), .vdd!(vdd!), .A(_681__20_), .Q(_465_) );
INX1 INX1_62 ( .gnd!(gnd!), .vdd!(vdd!), .A(PC1_20_), .Q(_466_) );
MU2IX1 MU2IX1_4 ( .gnd!(gnd!), .vdd!(vdd!), .IN0(_465_), .IN1(_466_), .Q(ALU_a_20_), .S(CTRL_IDEC1_cu_auipc_inst_bF_buf4) );
INX1 INX1_63 ( .gnd!(gnd!), .vdd!(vdd!), .A(_681__21_), .Q(_467_) );
INX1 INX1_64 ( .gnd!(gnd!), .vdd!(vdd!), .A(PC1_21_), .Q(_468_) );
MU2IX1 MU2IX1_5 ( .gnd!(gnd!), .vdd!(vdd!), .IN0(_467_), .IN1(_468_), .Q(ALU_a_21_), .S(CTRL_IDEC1_cu_auipc_inst_bF_buf4) );
MU2X1 MU2X1_39 ( .gnd!(gnd!), .vdd!(vdd!), .IN0(_681__22_), .IN1(PC1_22_), .Q(ALU_a_22_), .S(CTRL_IDEC1_cu_auipc_inst_bF_buf4) );
MU2X1 MU2X1_40 ( .gnd!(gnd!), .vdd!(vdd!), .IN0(_681__23_), .IN1(PC1_23_), .Q(ALU_a_23_), .S(CTRL_IDEC1_cu_auipc_inst_bF_buf2) );
MU2X1 MU2X1_41 ( .gnd!(gnd!), .vdd!(vdd!), .IN0(_681__24_), .IN1(PC1_24_), .Q(ALU_a_24_), .S(CTRL_IDEC1_cu_auipc_inst_bF_buf3) );
MU2X1 MU2X1_42 ( .gnd!(gnd!), .vdd!(vdd!), .IN0(_681__25_), .IN1(PC1_25_), .Q(ALU_a_25_), .S(CTRL_IDEC1_cu_auipc_inst_bF_buf3) );
MU2X1 MU2X1_43 ( .gnd!(gnd!), .vdd!(vdd!), .IN0(_681__26_), .IN1(PC1_26_), .Q(ALU_a_26_), .S(CTRL_IDEC1_cu_auipc_inst_bF_buf3) );
MU2X1 MU2X1_44 ( .gnd!(gnd!), .vdd!(vdd!), .IN0(_681__27_), .IN1(PC1_27_), .Q(ALU_a_27_), .S(CTRL_IDEC1_cu_auipc_inst_bF_buf2) );
INX1 INX1_65 ( .gnd!(gnd!), .vdd!(vdd!), .A(_681__28_), .Q(_469_) );
INX1 INX1_66 ( .gnd!(gnd!), .vdd!(vdd!), .A(PC1_28_), .Q(_470_) );
MU2IX1 MU2IX1_6 ( .gnd!(gnd!), .vdd!(vdd!), .IN0(_469_), .IN1(_470_), .Q(ALU_a_28_), .S(CTRL_IDEC1_cu_auipc_inst_bF_buf3) );
MU2X1 MU2X1_45 ( .gnd!(gnd!), .vdd!(vdd!), .IN0(_681__29_), .IN1(PC1_29_), .Q(ALU_a_29_), .S(CTRL_IDEC1_cu_auipc_inst_bF_buf2) );
MU2X1 MU2X1_46 ( .gnd!(gnd!), .vdd!(vdd!), .IN0(_681__30_), .IN1(PC1_30_), .Q(ALU_a_30_), .S(CTRL_IDEC1_cu_auipc_inst_bF_buf3) );
MU2X1 MU2X1_47 ( .gnd!(gnd!), .vdd!(vdd!), .IN0(_681__31_), .IN1(PC1_31_), .Q(ALU_a_31_), .S(CTRL_IDEC1_cu_auipc_inst_bF_buf3) );
MU2X1 MU2X1_48 ( .gnd!(gnd!), .vdd!(vdd!), .IN0(_678__0_), .IN1(I1_0_), .Q(ALU_b_0_), .S(CTRL_cu_alu_b_src_bF_buf0) );
MU2X1 MU2X1_49 ( .gnd!(gnd!), .vdd!(vdd!), .IN0(_678__1_), .IN1(I1_1_), .Q(ALU_b_1_), .S(CTRL_cu_alu_b_src_bF_buf1) );
MU2X1 MU2X1_50 ( .gnd!(gnd!), .vdd!(vdd!), .IN0(_678__2_), .IN1(I1_2_), .Q(ALU_b_2_), .S(CTRL_cu_alu_b_src_bF_buf3) );
MU2X1 MU2X1_51 ( .gnd!(gnd!), .vdd!(vdd!), .IN0(_678__3_), .IN1(I1_3_), .Q(ALU_b_3_), .S(CTRL_cu_alu_b_src_bF_buf3) );
MU2X1 MU2X1_52 ( .gnd!(gnd!), .vdd!(vdd!), .IN0(_678__4_), .IN1(I1_4_), .Q(ALU_b_4_), .S(CTRL_cu_alu_b_src_bF_buf3) );
MU2X1 MU2X1_53 ( .gnd!(gnd!), .vdd!(vdd!), .IN0(_678__5_), .IN1(I1_5_), .Q(ALU_b_5_), .S(CTRL_cu_alu_b_src_bF_buf3) );
MU2X1 MU2X1_54 ( .gnd!(gnd!), .vdd!(vdd!), .IN0(_678__6_), .IN1(I1_6_), .Q(ALU_b_6_), .S(CTRL_cu_alu_b_src_bF_buf3) );
MU2X1 MU2X1_55 ( .gnd!(gnd!), .vdd!(vdd!), .IN0(_678__7_), .IN1(I1_7_), .Q(ALU_b_7_), .S(CTRL_cu_alu_b_src_bF_buf4) );
MU2X1 MU2X1_56 ( .gnd!(gnd!), .vdd!(vdd!), .IN0(_678__8_), .IN1(I1_8_), .Q(ALU_b_8_), .S(CTRL_cu_alu_b_src_bF_buf3) );
MU2X1 MU2X1_57 ( .gnd!(gnd!), .vdd!(vdd!), .IN0(_678__9_), .IN1(I1_9_), .Q(ALU_b_9_), .S(CTRL_cu_alu_b_src_bF_buf3) );
MU2X1 MU2X1_58 ( .gnd!(gnd!), .vdd!(vdd!), .IN0(_678__10_), .IN1(I1_10_), .Q(ALU_b_10_), .S(CTRL_cu_alu_b_src_bF_buf4) );
MU2X1 MU2X1_59 ( .gnd!(gnd!), .vdd!(vdd!), .IN0(_678__11_), .IN1(I1_11_), .Q(ALU_b_11_), .S(CTRL_cu_alu_b_src_bF_buf4) );
MU2X1 MU2X1_60 ( .gnd!(gnd!), .vdd!(vdd!), .IN0(_678__12_), .IN1(I1_12_), .Q(ALU_b_12_), .S(CTRL_cu_alu_b_src_bF_buf4) );
MU2X1 MU2X1_61 ( .gnd!(gnd!), .vdd!(vdd!), .IN0(_678__13_), .IN1(I1_13_), .Q(ALU_b_13_), .S(CTRL_cu_alu_b_src_bF_buf4) );
MU2X1 MU2X1_62 ( .gnd!(gnd!), .vdd!(vdd!), .IN0(_678__14_), .IN1(I1_14_), .Q(ALU_b_14_), .S(CTRL_cu_alu_b_src_bF_buf4) );
MU2X1 MU2X1_63 ( .gnd!(gnd!), .vdd!(vdd!), .IN0(_678__15_), .IN1(I1_15_), .Q(ALU_b_15_), .S(CTRL_cu_alu_b_src_bF_buf4) );
MU2X1 MU2X1_64 ( .gnd!(gnd!), .vdd!(vdd!), .IN0(_678__16_), .IN1(I1_16_), .Q(ALU_b_16_), .S(CTRL_cu_alu_b_src_bF_buf1) );
MU2X1 MU2X1_65 ( .gnd!(gnd!), .vdd!(vdd!), .IN0(_678__17_), .IN1(I1_17_), .Q(ALU_b_17_), .S(CTRL_cu_alu_b_src_bF_buf0) );
MU2X1 MU2X1_66 ( .gnd!(gnd!), .vdd!(vdd!), .IN0(_678__18_), .IN1(I1_18_), .Q(ALU_b_18_), .S(CTRL_cu_alu_b_src_bF_buf1) );
MU2X1 MU2X1_67 ( .gnd!(gnd!), .vdd!(vdd!), .IN0(_678__19_), .IN1(I1_19_), .Q(ALU_b_19_), .S(CTRL_cu_alu_b_src_bF_buf0) );
MU2X1 MU2X1_68 ( .gnd!(gnd!), .vdd!(vdd!), .IN0(_678__20_), .IN1(I1_20_), .Q(ALU_b_20_), .S(CTRL_cu_alu_b_src_bF_buf2) );
MU2X1 MU2X1_69 ( .gnd!(gnd!), .vdd!(vdd!), .IN0(_678__21_), .IN1(I1_21_), .Q(ALU_b_21_), .S(CTRL_cu_alu_b_src_bF_buf1) );
MU2X1 MU2X1_70 ( .gnd!(gnd!), .vdd!(vdd!), .IN0(_678__22_), .IN1(I1_22_), .Q(ALU_b_22_), .S(CTRL_cu_alu_b_src_bF_buf0) );
MU2X1 MU2X1_71 ( .gnd!(gnd!), .vdd!(vdd!), .IN0(_678__23_), .IN1(I1_23_), .Q(ALU_b_23_), .S(CTRL_cu_alu_b_src_bF_buf0) );
MU2X1 MU2X1_72 ( .gnd!(gnd!), .vdd!(vdd!), .IN0(_678__24_), .IN1(I1_24_), .Q(ALU_b_24_), .S(CTRL_cu_alu_b_src_bF_buf2) );
MU2X1 MU2X1_73 ( .gnd!(gnd!), .vdd!(vdd!), .IN0(_678__25_), .IN1(I1_25_), .Q(ALU_b_25_), .S(CTRL_cu_alu_b_src_bF_buf2) );
MU2X1 MU2X1_74 ( .gnd!(gnd!), .vdd!(vdd!), .IN0(_678__26_), .IN1(I1_26_), .Q(ALU_b_26_), .S(CTRL_cu_alu_b_src_bF_buf2) );
MU2X1 MU2X1_75 ( .gnd!(gnd!), .vdd!(vdd!), .IN0(_678__27_), .IN1(I1_27_), .Q(ALU_b_27_), .S(CTRL_cu_alu_b_src_bF_buf1) );
MU2X1 MU2X1_76 ( .gnd!(gnd!), .vdd!(vdd!), .IN0(_678__28_), .IN1(I1_28_), .Q(ALU_b_28_), .S(CTRL_cu_alu_b_src_bF_buf1) );
MU2X1 MU2X1_77 ( .gnd!(gnd!), .vdd!(vdd!), .IN0(_678__29_), .IN1(I1_29_), .Q(ALU_b_29_), .S(CTRL_cu_alu_b_src_bF_buf0) );
MU2X1 MU2X1_78 ( .gnd!(gnd!), .vdd!(vdd!), .IN0(_678__30_), .IN1(I1_30_), .Q(ALU_b_30_), .S(CTRL_cu_alu_b_src_bF_buf2) );
MU2X1 MU2X1_79 ( .gnd!(gnd!), .vdd!(vdd!), .IN0(_678__31_), .IN1(I1_31_), .Q(ALU_b_31_), .S(CTRL_cu_alu_b_src_bF_buf2) );
ON21X1 ON21X1_128 ( .gnd!(gnd!), .vdd!(vdd!), .A(_28_), .B(CTRL_cyc_bF_buf2_bF_buf0), .C(_593_), .Q(_677__0_) );
ON21X1 ON21X1_129 ( .gnd!(gnd!), .vdd!(vdd!), .A(_46_), .B(CTRL_cyc_bF_buf1_bF_buf2), .C(_597_), .Q(_677__1_) );
ON21X1 ON21X1_130 ( .gnd!(gnd!), .vdd!(vdd!), .A(_59_), .B(CTRL_cyc_bF_buf0_bF_buf3), .C(_600_), .Q(_677__2_) );
ON21X1 ON21X1_131 ( .gnd!(gnd!), .vdd!(vdd!), .A(_71_), .B(CTRL_cyc_bF_buf14_bF_buf1), .C(_603_), .Q(_677__3_) );
ON21X1 ON21X1_132 ( .gnd!(gnd!), .vdd!(vdd!), .A(_84_), .B(CTRL_cyc_bF_buf13_bF_buf1), .C(_606_), .Q(_677__4_) );
ON21X1 ON21X1_133 ( .gnd!(gnd!), .vdd!(vdd!), .A(_96_), .B(CTRL_cyc_bF_buf12_bF_buf1), .C(_609_), .Q(_677__5_) );
ON21X1 ON21X1_134 ( .gnd!(gnd!), .vdd!(vdd!), .A(_109_), .B(CTRL_cyc_bF_buf11_bF_buf0), .C(_612_), .Q(_677__6_) );
ON21X1 ON21X1_135 ( .gnd!(gnd!), .vdd!(vdd!), .A(_121_), .B(CTRL_cyc_bF_buf10_bF_buf3), .C(_615_), .Q(_677__7_) );
ON21X1 ON21X1_136 ( .gnd!(gnd!), .vdd!(vdd!), .A(_133_), .B(CTRL_cyc_bF_buf9_bF_buf0), .C(_618_), .Q(_677__8_) );
ON21X1 ON21X1_137 ( .gnd!(gnd!), .vdd!(vdd!), .A(_146_), .B(CTRL_cyc_bF_buf8_bF_buf2), .C(_621_), .Q(_677__9_) );
ON21X1 ON21X1_138 ( .gnd!(gnd!), .vdd!(vdd!), .A(_159_), .B(CTRL_cyc_bF_buf7_bF_buf3), .C(_624_), .Q(_677__10_) );
ON21X1 ON21X1_139 ( .gnd!(gnd!), .vdd!(vdd!), .A(_172_), .B(CTRL_cyc_bF_buf6_bF_buf0), .C(_627_), .Q(_677__11_) );
ON21X1 ON21X1_140 ( .gnd!(gnd!), .vdd!(vdd!), .A(_185_), .B(CTRL_cyc_bF_buf5_bF_buf2), .C(_630_), .Q(_677__12_) );
ON21X1 ON21X1_141 ( .gnd!(gnd!), .vdd!(vdd!), .A(_197_), .B(CTRL_cyc_bF_buf4_bF_buf3), .C(_633_), .Q(_677__13_) );
ON21X1 ON21X1_142 ( .gnd!(gnd!), .vdd!(vdd!), .A(_210_), .B(CTRL_cyc_bF_buf3_bF_buf3), .C(_636_), .Q(_677__14_) );
ON21X1 ON21X1_143 ( .gnd!(gnd!), .vdd!(vdd!), .A(_223_), .B(CTRL_cyc_bF_buf2_bF_buf0), .C(_639_), .Q(_677__15_) );
ON21X1 ON21X1_144 ( .gnd!(gnd!), .vdd!(vdd!), .A(_235_), .B(CTRL_cyc_bF_buf1_bF_buf3), .C(_642_), .Q(_677__16_) );
ON21X1 ON21X1_145 ( .gnd!(gnd!), .vdd!(vdd!), .A(_248_), .B(CTRL_cyc_bF_buf0_bF_buf2), .C(_645_), .Q(_677__17_) );
ON21X1 ON21X1_146 ( .gnd!(gnd!), .vdd!(vdd!), .A(_261_), .B(CTRL_cyc_bF_buf14_bF_buf0), .C(_648_), .Q(_677__18_) );
ON21X1 ON21X1_147 ( .gnd!(gnd!), .vdd!(vdd!), .A(_275_), .B(CTRL_cyc_bF_buf13_bF_buf1), .C(_651_), .Q(_677__19_) );
ON21X1 ON21X1_148 ( .gnd!(gnd!), .vdd!(vdd!), .A(_287_), .B(CTRL_cyc_bF_buf12_bF_buf1), .C(_654_), .Q(_677__20_) );
ON21X1 ON21X1_149 ( .gnd!(gnd!), .vdd!(vdd!), .A(_299_), .B(CTRL_cyc_bF_buf11_bF_buf2), .C(_657_), .Q(_677__21_) );
ON21X1 ON21X1_150 ( .gnd!(gnd!), .vdd!(vdd!), .A(_312_), .B(CTRL_cyc_bF_buf10_bF_buf3), .C(_660_), .Q(_677__22_) );
ON21X1 ON21X1_151 ( .gnd!(gnd!), .vdd!(vdd!), .A(_325_), .B(CTRL_cyc_bF_buf9_bF_buf3), .C(_663_), .Q(_677__23_) );
ON21X1 ON21X1_152 ( .gnd!(gnd!), .vdd!(vdd!), .A(_338_), .B(CTRL_cyc_bF_buf8_bF_buf2), .C(_666_), .Q(_677__24_) );
ON21X1 ON21X1_153 ( .gnd!(gnd!), .vdd!(vdd!), .A(_351_), .B(CTRL_cyc_bF_buf7_bF_buf1), .C(_669_), .Q(_677__25_) );
ON21X1 ON21X1_154 ( .gnd!(gnd!), .vdd!(vdd!), .A(_364_), .B(CTRL_cyc_bF_buf6_bF_buf2), .C(_672_), .Q(_677__26_) );
ON21X1 ON21X1_155 ( .gnd!(gnd!), .vdd!(vdd!), .A(_376_), .B(CTRL_cyc_bF_buf5_bF_buf1), .C(_675_), .Q(_677__27_) );
ON21X1 ON21X1_156 ( .gnd!(gnd!), .vdd!(vdd!), .A(_388_), .B(CTRL_cyc_bF_buf4_bF_buf0), .C(_8_), .Q(_677__28_) );
ON21X1 ON21X1_157 ( .gnd!(gnd!), .vdd!(vdd!), .A(_401_), .B(CTRL_cyc_bF_buf3_bF_buf3), .C(_11_), .Q(_677__29_) );
ON21X1 ON21X1_158 ( .gnd!(gnd!), .vdd!(vdd!), .A(_414_), .B(CTRL_cyc_bF_buf2_bF_buf1), .C(_14_), .Q(_677__30_) );
ON21X1 ON21X1_159 ( .gnd!(gnd!), .vdd!(vdd!), .A(_427_), .B(CTRL_cyc_bF_buf1_bF_buf0), .C(_17_), .Q(_677__31_) );
AND2X2 AND2X2_1 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_cyc_bF_buf0_bF_buf0), .B(_682__0_bF_buf3), .Q(_679__0_) );
NA2I1X1 NA2I1X1_33 ( .gnd!(gnd!), .vdd!(vdd!), .AN(_682__1_bF_buf4), .B(CTRL_cyc_bF_buf14_bF_buf2), .Q(_679__1_) );
INX3 INX3_4 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_cu_r1_ld), .Q(_471_) );
NA2X1 NA2X1_99 ( .gnd!(gnd!), .vdd!(vdd!), .A(_471__bF_buf2), .B(_681__0_), .Q(_472_) );
INX3 INX3_5 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_cu_r1_src_bF_buf2), .Q(_473_) );
NO2X1 NO2X1_89 ( .gnd!(gnd!), .vdd!(vdd!), .A(_686__1_), .B(_686__0_), .Q(_474_) );
NO2X1 NO2X1_90 ( .gnd!(gnd!), .vdd!(vdd!), .A(_686__3_), .B(_686__2_), .Q(_475_) );
NA3I1X2 NA3I1X2_2 ( .gnd!(gnd!), .vdd!(vdd!), .AN(_686__4_), .B(_474_), .C(_475_), .Q(_476_) );
NA2X1 NA2X1_100 ( .gnd!(gnd!), .vdd!(vdd!), .A(_476__bF_buf3), .B(rfRS1[0]), .Q(_477_) );
AN21X1 AN21X1_45 ( .gnd!(gnd!), .vdd!(vdd!), .A(_477_), .B(_473__bF_buf4), .C(_471__bF_buf4), .Q(_478_) );
ON21X1 ON21X1_160 ( .gnd!(gnd!), .vdd!(vdd!), .A(_34_), .B(_473__bF_buf3), .C(_478_), .Q(_479_) );
NA2X1 NA2X1_101 ( .gnd!(gnd!), .vdd!(vdd!), .A(_479_), .B(_472_), .Q(_3__0_) );
ON211X1 ON211X1_23 ( .gnd!(gnd!), .vdd!(vdd!), .A(_48_), .B(_49_), .C(CTRL_cu_r1_src_bF_buf3), .D(_41_), .Q(_480_) );
AN21X1 AN21X1_46 ( .gnd!(gnd!), .vdd!(vdd!), .A(_476__bF_buf1), .B(rfRS1[1]), .C(CTRL_cu_r1_src_bF_buf1), .Q(_481_) );
NO2X1 NO2X1_91 ( .gnd!(gnd!), .vdd!(vdd!), .A(_471__bF_buf1), .B(_481_), .Q(_482_) );
AO22X2 AO22X2_12 ( .gnd!(gnd!), .vdd!(vdd!), .A(_681__1_), .B(_471__bF_buf2), .C(_480_), .D(_482_), .Q(_3__1_) );
NA2X1 NA2X1_102 ( .gnd!(gnd!), .vdd!(vdd!), .A(_471__bF_buf2), .B(_681__2_), .Q(_483_) );
NA2X1 NA2X1_103 ( .gnd!(gnd!), .vdd!(vdd!), .A(_476__bF_buf2), .B(rfRS1[2]), .Q(_484_) );
AN21X1 AN21X1_47 ( .gnd!(gnd!), .vdd!(vdd!), .A(_484_), .B(_473__bF_buf5), .C(_471__bF_buf0), .Q(_485_) );
ON21X1 ON21X1_161 ( .gnd!(gnd!), .vdd!(vdd!), .A(_63_), .B(_473__bF_buf1), .C(_485_), .Q(_486_) );
NA2X1 NA2X1_104 ( .gnd!(gnd!), .vdd!(vdd!), .A(_486_), .B(_483_), .Q(_3__2_) );
ON211X1 ON211X1_24 ( .gnd!(gnd!), .vdd!(vdd!), .A(_73_), .B(_74_), .C(CTRL_cu_r1_src_bF_buf3), .D(_66_), .Q(_487_) );
AN21X1 AN21X1_48 ( .gnd!(gnd!), .vdd!(vdd!), .A(_476__bF_buf3), .B(rfRS1[3]), .C(CTRL_cu_r1_src_bF_buf2), .Q(_488_) );
NO2X1 NO2X1_92 ( .gnd!(gnd!), .vdd!(vdd!), .A(_471__bF_buf4), .B(_488_), .Q(_489_) );
AO22X2 AO22X2_13 ( .gnd!(gnd!), .vdd!(vdd!), .A(_681__3_), .B(_471__bF_buf2), .C(_487_), .D(_489_), .Q(_3__3_) );
NA2X1 NA2X1_105 ( .gnd!(gnd!), .vdd!(vdd!), .A(_471__bF_buf7), .B(_681__4_), .Q(_490_) );
NA2X1 NA2X1_106 ( .gnd!(gnd!), .vdd!(vdd!), .A(_476__bF_buf2), .B(rfRS1[4]), .Q(_491_) );
AN21X1 AN21X1_49 ( .gnd!(gnd!), .vdd!(vdd!), .A(_491_), .B(_473__bF_buf5), .C(_471__bF_buf0), .Q(_492_) );
ON21X1 ON21X1_162 ( .gnd!(gnd!), .vdd!(vdd!), .A(_88_), .B(_473__bF_buf1), .C(_492_), .Q(_493_) );
NA2X1 NA2X1_107 ( .gnd!(gnd!), .vdd!(vdd!), .A(_493_), .B(_490_), .Q(_3__4_) );
ON211X1 ON211X1_25 ( .gnd!(gnd!), .vdd!(vdd!), .A(_98_), .B(_99_), .C(CTRL_cu_r1_src_bF_buf3), .D(_91_), .Q(_494_) );
NA2X1 NA2X1_108 ( .gnd!(gnd!), .vdd!(vdd!), .A(_476__bF_buf3), .B(rfRS1[5]), .Q(_495_) );
AN21X1 AN21X1_50 ( .gnd!(gnd!), .vdd!(vdd!), .A(_495_), .B(_473__bF_buf4), .C(_471__bF_buf4), .Q(_496_) );
AO22X2 AO22X2_14 ( .gnd!(gnd!), .vdd!(vdd!), .A(_681__5_), .B(_471__bF_buf2), .C(_494_), .D(_496_), .Q(_3__5_) );
NA2X1 NA2X1_109 ( .gnd!(gnd!), .vdd!(vdd!), .A(_471__bF_buf2), .B(_681__6_), .Q(_497_) );
NA2X1 NA2X1_110 ( .gnd!(gnd!), .vdd!(vdd!), .A(_476__bF_buf1), .B(rfRS1[6]), .Q(_498_) );
AN21X1 AN21X1_51 ( .gnd!(gnd!), .vdd!(vdd!), .A(_498_), .B(_473__bF_buf1), .C(_471__bF_buf1), .Q(_499_) );
ON21X1 ON21X1_163 ( .gnd!(gnd!), .vdd!(vdd!), .A(_113_), .B(_473__bF_buf1), .C(_499_), .Q(_500_) );
NA2X1 NA2X1_111 ( .gnd!(gnd!), .vdd!(vdd!), .A(_500_), .B(_497_), .Q(_3__6_) );
ON211X1 ON211X1_26 ( .gnd!(gnd!), .vdd!(vdd!), .A(_123_), .B(_124_), .C(CTRL_cu_r1_src_bF_buf0), .D(_116_), .Q(_501_) );
AN21X1 AN21X1_52 ( .gnd!(gnd!), .vdd!(vdd!), .A(_476__bF_buf0), .B(rfRS1[7]), .C(CTRL_cu_r1_src_bF_buf2), .Q(_502_) );
NO2X1 NO2X1_93 ( .gnd!(gnd!), .vdd!(vdd!), .A(_471__bF_buf7), .B(_502_), .Q(_503_) );
AO22X2 AO22X2_15 ( .gnd!(gnd!), .vdd!(vdd!), .A(_681__7_), .B(_471__bF_buf7), .C(_501_), .D(_503_), .Q(_3__7_) );
ON211X1 ON211X1_27 ( .gnd!(gnd!), .vdd!(vdd!), .A(_135_), .B(_136_), .C(CTRL_cu_r1_src_bF_buf0), .D(_128_), .Q(_504_) );
NA2X1 NA2X1_112 ( .gnd!(gnd!), .vdd!(vdd!), .A(_476__bF_buf1), .B(rfRS1[8]), .Q(_505_) );
AN21X1 AN21X1_53 ( .gnd!(gnd!), .vdd!(vdd!), .A(_505_), .B(_473__bF_buf1), .C(_471__bF_buf5), .Q(_506_) );
AO22X2 AO22X2_16 ( .gnd!(gnd!), .vdd!(vdd!), .A(_681__8_), .B(_471__bF_buf2), .C(_504_), .D(_506_), .Q(_3__8_) );
NA2X1 NA2X1_113 ( .gnd!(gnd!), .vdd!(vdd!), .A(_471__bF_buf6), .B(_681__9_), .Q(_507_) );
NA2X1 NA2X1_114 ( .gnd!(gnd!), .vdd!(vdd!), .A(_476__bF_buf0), .B(rfRS1[9]), .Q(_508_) );
AN21X1 AN21X1_54 ( .gnd!(gnd!), .vdd!(vdd!), .A(_508_), .B(_473__bF_buf5), .C(_471__bF_buf6), .Q(_509_) );
ON21X1 ON21X1_164 ( .gnd!(gnd!), .vdd!(vdd!), .A(_150_), .B(_473__bF_buf0), .C(_509_), .Q(_510_) );
NA2X1 NA2X1_115 ( .gnd!(gnd!), .vdd!(vdd!), .A(_510_), .B(_507_), .Q(_3__9_) );
NA2X1 NA2X1_116 ( .gnd!(gnd!), .vdd!(vdd!), .A(_471__bF_buf3), .B(_681__10_), .Q(_511_) );
NA2X1 NA2X1_117 ( .gnd!(gnd!), .vdd!(vdd!), .A(_476__bF_buf4), .B(rfRS1[10]), .Q(_512_) );
AN21X1 AN21X1_55 ( .gnd!(gnd!), .vdd!(vdd!), .A(_512_), .B(_473__bF_buf2), .C(_471__bF_buf3), .Q(_513_) );
ON21X1 ON21X1_165 ( .gnd!(gnd!), .vdd!(vdd!), .A(_163_), .B(_473__bF_buf2), .C(_513_), .Q(_514_) );
NA2X1 NA2X1_118 ( .gnd!(gnd!), .vdd!(vdd!), .A(_514_), .B(_511_), .Q(_3__10_) );
NA2X1 NA2X1_119 ( .gnd!(gnd!), .vdd!(vdd!), .A(_471__bF_buf2), .B(_681__11_), .Q(_515_) );
NA2X1 NA2X1_120 ( .gnd!(gnd!), .vdd!(vdd!), .A(_476__bF_buf3), .B(rfRS1[11]), .Q(_516_) );
AN21X1 AN21X1_56 ( .gnd!(gnd!), .vdd!(vdd!), .A(_516_), .B(_473__bF_buf4), .C(_471__bF_buf0), .Q(_517_) );
ON21X1 ON21X1_166 ( .gnd!(gnd!), .vdd!(vdd!), .A(_176_), .B(_473__bF_buf3), .C(_517_), .Q(_518_) );
NA2X1 NA2X1_121 ( .gnd!(gnd!), .vdd!(vdd!), .A(_518_), .B(_515_), .Q(_3__11_) );
NA2X1 NA2X1_122 ( .gnd!(gnd!), .vdd!(vdd!), .A(_471__bF_buf4), .B(_681__12_), .Q(_519_) );
NA2X1 NA2X1_123 ( .gnd!(gnd!), .vdd!(vdd!), .A(_476__bF_buf2), .B(rfRS1[12]), .Q(_520_) );
AN21X1 AN21X1_57 ( .gnd!(gnd!), .vdd!(vdd!), .A(_520_), .B(_473__bF_buf5), .C(_471__bF_buf0), .Q(_521_) );
ON21X1 ON21X1_167 ( .gnd!(gnd!), .vdd!(vdd!), .A(_189_), .B(_473__bF_buf4), .C(_521_), .Q(_522_) );
NA2X1 NA2X1_124 ( .gnd!(gnd!), .vdd!(vdd!), .A(_522_), .B(_519_), .Q(_3__12_) );
ON211X1 ON211X1_28 ( .gnd!(gnd!), .vdd!(vdd!), .A(_199_), .B(_200_), .C(CTRL_cu_r1_src_bF_buf0), .D(_192_), .Q(_523_) );
AN21X1 AN21X1_58 ( .gnd!(gnd!), .vdd!(vdd!), .A(_476__bF_buf0), .B(rfRS1[13]), .C(CTRL_cu_r1_src_bF_buf2), .Q(_524_) );
NO2X1 NO2X1_94 ( .gnd!(gnd!), .vdd!(vdd!), .A(_471__bF_buf5), .B(_524_), .Q(_525_) );
AO22X2 AO22X2_17 ( .gnd!(gnd!), .vdd!(vdd!), .A(_681__13_), .B(_471__bF_buf7), .C(_523_), .D(_525_), .Q(_3__13_) );
NA2X1 NA2X1_125 ( .gnd!(gnd!), .vdd!(vdd!), .A(_471__bF_buf1), .B(_681__14_), .Q(_526_) );
NA2X1 NA2X1_126 ( .gnd!(gnd!), .vdd!(vdd!), .A(_476__bF_buf3), .B(rfRS1[14]), .Q(_527_) );
AN21X1 AN21X1_59 ( .gnd!(gnd!), .vdd!(vdd!), .A(_527_), .B(_473__bF_buf3), .C(_471__bF_buf4), .Q(_528_) );
ON21X1 ON21X1_168 ( .gnd!(gnd!), .vdd!(vdd!), .A(_214_), .B(_473__bF_buf3), .C(_528_), .Q(_529_) );
NA2X1 NA2X1_127 ( .gnd!(gnd!), .vdd!(vdd!), .A(_529_), .B(_526_), .Q(_3__14_) );
NA2X1 NA2X1_128 ( .gnd!(gnd!), .vdd!(vdd!), .A(_471__bF_buf6), .B(_681__15_), .Q(_530_) );
NA2X1 NA2X1_129 ( .gnd!(gnd!), .vdd!(vdd!), .A(_476__bF_buf4), .B(rfRS1[15]), .Q(_531_) );
AN21X1 AN21X1_60 ( .gnd!(gnd!), .vdd!(vdd!), .A(_531_), .B(_473__bF_buf0), .C(_471__bF_buf6), .Q(_532_) );
ON21X1 ON21X1_169 ( .gnd!(gnd!), .vdd!(vdd!), .A(_227_), .B(_473__bF_buf0), .C(_532_), .Q(_533_) );
NA2X1 NA2X1_130 ( .gnd!(gnd!), .vdd!(vdd!), .A(_533_), .B(_530_), .Q(_3__15_) );
ON211X1 ON211X1_29 ( .gnd!(gnd!), .vdd!(vdd!), .A(_237_), .B(_238_), .C(CTRL_cu_r1_src_bF_buf1), .D(_230_), .Q(_534_) );
NA2X1 NA2X1_131 ( .gnd!(gnd!), .vdd!(vdd!), .A(_476__bF_buf1), .B(rfRS1[16]), .Q(_535_) );
AN21X1 AN21X1_61 ( .gnd!(gnd!), .vdd!(vdd!), .A(_535_), .B(_473__bF_buf1), .C(_471__bF_buf5), .Q(_536_) );
AO22X2 AO22X2_18 ( .gnd!(gnd!), .vdd!(vdd!), .A(_681__16_), .B(_471__bF_buf7), .C(_534_), .D(_536_), .Q(_3__16_) );
NA2X1 NA2X1_132 ( .gnd!(gnd!), .vdd!(vdd!), .A(_471__bF_buf5), .B(_681__17_), .Q(_537_) );
NA2X1 NA2X1_133 ( .gnd!(gnd!), .vdd!(vdd!), .A(_476__bF_buf0), .B(rfRS1[17]), .Q(_538_) );
AN21X1 AN21X1_62 ( .gnd!(gnd!), .vdd!(vdd!), .A(_538_), .B(_473__bF_buf5), .C(_471__bF_buf0), .Q(_539_) );
ON21X1 ON21X1_170 ( .gnd!(gnd!), .vdd!(vdd!), .A(_252_), .B(_473__bF_buf4), .C(_539_), .Q(_540_) );
NA2X1 NA2X1_134 ( .gnd!(gnd!), .vdd!(vdd!), .A(_540_), .B(_537_), .Q(_3__17_) );
NA2X1 NA2X1_135 ( .gnd!(gnd!), .vdd!(vdd!), .A(_471__bF_buf1), .B(_681__18_), .Q(_541_) );
NA2X1 NA2X1_136 ( .gnd!(gnd!), .vdd!(vdd!), .A(_476__bF_buf3), .B(rfRS1[18]), .Q(_542_) );
AN21X1 AN21X1_63 ( .gnd!(gnd!), .vdd!(vdd!), .A(_542_), .B(_473__bF_buf3), .C(_471__bF_buf4), .Q(_543_) );
ON21X1 ON21X1_171 ( .gnd!(gnd!), .vdd!(vdd!), .A(_265_), .B(_473__bF_buf3), .C(_543_), .Q(_544_) );
NA2X1 NA2X1_137 ( .gnd!(gnd!), .vdd!(vdd!), .A(_544_), .B(_541_), .Q(_3__18_) );
NA2X1 NA2X1_138 ( .gnd!(gnd!), .vdd!(vdd!), .A(_471__bF_buf3), .B(_681__19_), .Q(_545_) );
NA2X1 NA2X1_139 ( .gnd!(gnd!), .vdd!(vdd!), .A(_476__bF_buf4), .B(rfRS1[19]), .Q(_546_) );
AN21X1 AN21X1_64 ( .gnd!(gnd!), .vdd!(vdd!), .A(_546_), .B(_473__bF_buf2), .C(_471__bF_buf3), .Q(_547_) );
ON21X1 ON21X1_172 ( .gnd!(gnd!), .vdd!(vdd!), .A(_279_), .B(_473__bF_buf2), .C(_547_), .Q(_548_) );
NA2X1 NA2X1_140 ( .gnd!(gnd!), .vdd!(vdd!), .A(_548_), .B(_545_), .Q(_3__19_) );
ON211X1 ON211X1_30 ( .gnd!(gnd!), .vdd!(vdd!), .A(_289_), .B(_290_), .C(CTRL_cu_r1_src_bF_buf0), .D(_282_), .Q(_549_) );
NA2X1 NA2X1_141 ( .gnd!(gnd!), .vdd!(vdd!), .A(_476__bF_buf2), .B(rfRS1[20]), .Q(_550_) );
AN21X1 AN21X1_65 ( .gnd!(gnd!), .vdd!(vdd!), .A(_550_), .B(_473__bF_buf1), .C(_471__bF_buf1), .Q(_551_) );
AO22X2 AO22X2_19 ( .gnd!(gnd!), .vdd!(vdd!), .A(_681__20_), .B(_471__bF_buf7), .C(_549_), .D(_551_), .Q(_3__20_) );
ON211X1 ON211X1_31 ( .gnd!(gnd!), .vdd!(vdd!), .A(_301_), .B(_302_), .C(CTRL_cu_r1_src_bF_buf3), .D(_294_), .Q(_552_) );
NA2X1 NA2X1_142 ( .gnd!(gnd!), .vdd!(vdd!), .A(_476__bF_buf0), .B(rfRS1[21]), .Q(_553_) );
AN21X1 AN21X1_66 ( .gnd!(gnd!), .vdd!(vdd!), .A(_553_), .B(_473__bF_buf0), .C(_471__bF_buf5), .Q(_554_) );
AO22X2 AO22X2_20 ( .gnd!(gnd!), .vdd!(vdd!), .A(_681__21_), .B(_471__bF_buf7), .C(_552_), .D(_554_), .Q(_3__21_) );
NA2X1 NA2X1_143 ( .gnd!(gnd!), .vdd!(vdd!), .A(_471__bF_buf3), .B(_681__22_), .Q(_555_) );
NA2X1 NA2X1_144 ( .gnd!(gnd!), .vdd!(vdd!), .A(_476__bF_buf4), .B(rfRS1[22]), .Q(_556_) );
AN21X1 AN21X1_67 ( .gnd!(gnd!), .vdd!(vdd!), .A(_556_), .B(_473__bF_buf2), .C(_471__bF_buf3), .Q(_557_) );
ON21X1 ON21X1_173 ( .gnd!(gnd!), .vdd!(vdd!), .A(_316_), .B(_473__bF_buf2), .C(_557_), .Q(_558_) );
NA2X1 NA2X1_145 ( .gnd!(gnd!), .vdd!(vdd!), .A(_558_), .B(_555_), .Q(_3__22_) );
NA2X1 NA2X1_146 ( .gnd!(gnd!), .vdd!(vdd!), .A(_471__bF_buf4), .B(_681__23_), .Q(_559_) );
NA2X1 NA2X1_147 ( .gnd!(gnd!), .vdd!(vdd!), .A(_476__bF_buf2), .B(rfRS1[23]), .Q(_560_) );
AN21X1 AN21X1_68 ( .gnd!(gnd!), .vdd!(vdd!), .A(_560_), .B(_473__bF_buf4), .C(_471__bF_buf0), .Q(_561_) );
ON21X1 ON21X1_174 ( .gnd!(gnd!), .vdd!(vdd!), .A(_329_), .B(_473__bF_buf4), .C(_561_), .Q(_562_) );
NA2X1 NA2X1_148 ( .gnd!(gnd!), .vdd!(vdd!), .A(_562_), .B(_559_), .Q(_3__23_) );
NA2X1 NA2X1_149 ( .gnd!(gnd!), .vdd!(vdd!), .A(_471__bF_buf6), .B(_681__24_), .Q(_563_) );
NA2X1 NA2X1_150 ( .gnd!(gnd!), .vdd!(vdd!), .A(_476__bF_buf0), .B(rfRS1[24]), .Q(_564_) );
AN21X1 AN21X1_69 ( .gnd!(gnd!), .vdd!(vdd!), .A(_564_), .B(_473__bF_buf5), .C(_471__bF_buf6), .Q(_565_) );
ON21X1 ON21X1_175 ( .gnd!(gnd!), .vdd!(vdd!), .A(_342_), .B(_473__bF_buf5), .C(_565_), .Q(_566_) );
NA2X1 NA2X1_151 ( .gnd!(gnd!), .vdd!(vdd!), .A(_566_), .B(_563_), .Q(_3__24_) );
NA2X1 NA2X1_152 ( .gnd!(gnd!), .vdd!(vdd!), .A(_471__bF_buf1), .B(_681__25_), .Q(_567_) );
NA2X1 NA2X1_153 ( .gnd!(gnd!), .vdd!(vdd!), .A(_476__bF_buf3), .B(rfRS1[25]), .Q(_568_) );
AN21X1 AN21X1_70 ( .gnd!(gnd!), .vdd!(vdd!), .A(_568_), .B(_473__bF_buf3), .C(_471__bF_buf4), .Q(_569_) );
ON21X1 ON21X1_176 ( .gnd!(gnd!), .vdd!(vdd!), .A(_355_), .B(_473__bF_buf3), .C(_569_), .Q(_570_) );
NA2X1 NA2X1_154 ( .gnd!(gnd!), .vdd!(vdd!), .A(_570_), .B(_567_), .Q(_3__25_) );
NA2X1 NA2X1_155 ( .gnd!(gnd!), .vdd!(vdd!), .A(_471__bF_buf0), .B(_681__26_), .Q(_571_) );
NA2X1 NA2X1_156 ( .gnd!(gnd!), .vdd!(vdd!), .A(_476__bF_buf2), .B(rfRS1[26]), .Q(_572_) );
AN21X1 AN21X1_71 ( .gnd!(gnd!), .vdd!(vdd!), .A(_572_), .B(_473__bF_buf5), .C(_471__bF_buf0), .Q(_573_) );
ON21X1 ON21X1_177 ( .gnd!(gnd!), .vdd!(vdd!), .A(_368_), .B(_473__bF_buf4), .C(_573_), .Q(_574_) );
NA2X1 NA2X1_157 ( .gnd!(gnd!), .vdd!(vdd!), .A(_574_), .B(_571_), .Q(_3__26_) );
ON211X1 ON211X1_32 ( .gnd!(gnd!), .vdd!(vdd!), .A(_378_), .B(_379_), .C(CTRL_cu_r1_src_bF_buf1), .D(_371_), .Q(_575_) );
AN21X1 AN21X1_72 ( .gnd!(gnd!), .vdd!(vdd!), .A(_476__bF_buf1), .B(rfRS1[27]), .C(CTRL_cu_r1_src_bF_buf1), .Q(_576_) );
NO2X1 NO2X1_95 ( .gnd!(gnd!), .vdd!(vdd!), .A(_471__bF_buf5), .B(_576_), .Q(_577_) );
AO22X2 AO22X2_21 ( .gnd!(gnd!), .vdd!(vdd!), .A(_681__27_), .B(_471__bF_buf7), .C(_575_), .D(_577_), .Q(_3__27_) );
ON211X1 ON211X1_33 ( .gnd!(gnd!), .vdd!(vdd!), .A(_390_), .B(_391_), .C(CTRL_cu_r1_src_bF_buf3), .D(_383_), .Q(_578_) );
NA2X1 NA2X1_158 ( .gnd!(gnd!), .vdd!(vdd!), .A(_476__bF_buf1), .B(rfRS1[28]), .Q(_579_) );
AN21X1 AN21X1_73 ( .gnd!(gnd!), .vdd!(vdd!), .A(_579_), .B(_473__bF_buf1), .C(_471__bF_buf1), .Q(_580_) );
AO22X2 AO22X2_22 ( .gnd!(gnd!), .vdd!(vdd!), .A(_681__28_), .B(_471__bF_buf1), .C(_578_), .D(_580_), .Q(_3__28_) );
NA2X1 NA2X1_159 ( .gnd!(gnd!), .vdd!(vdd!), .A(_471__bF_buf5), .B(_681__29_), .Q(_581_) );
NA2X1 NA2X1_160 ( .gnd!(gnd!), .vdd!(vdd!), .A(_476__bF_buf4), .B(rfRS1[29]), .Q(_582_) );
AN21X1 AN21X1_74 ( .gnd!(gnd!), .vdd!(vdd!), .A(_582_), .B(_473__bF_buf0), .C(_471__bF_buf6), .Q(_583_) );
ON21X1 ON21X1_178 ( .gnd!(gnd!), .vdd!(vdd!), .A(_405_), .B(_473__bF_buf0), .C(_583_), .Q(_584_) );
NA2X1 NA2X1_161 ( .gnd!(gnd!), .vdd!(vdd!), .A(_584_), .B(_581_), .Q(_3__29_) );
NA2X1 NA2X1_162 ( .gnd!(gnd!), .vdd!(vdd!), .A(_471__bF_buf3), .B(_681__30_), .Q(_585_) );
NA2X1 NA2X1_163 ( .gnd!(gnd!), .vdd!(vdd!), .A(_476__bF_buf4), .B(rfRS1[30]), .Q(_586_) );
AN21X1 AN21X1_75 ( .gnd!(gnd!), .vdd!(vdd!), .A(_586_), .B(_473__bF_buf2), .C(_471__bF_buf3), .Q(_587_) );
ON21X1 ON21X1_179 ( .gnd!(gnd!), .vdd!(vdd!), .A(_418_), .B(_473__bF_buf2), .C(_587_), .Q(_588_) );
NA2X1 NA2X1_164 ( .gnd!(gnd!), .vdd!(vdd!), .A(_588_), .B(_585_), .Q(_3__30_) );
NA2X1 NA2X1_165 ( .gnd!(gnd!), .vdd!(vdd!), .A(_471__bF_buf5), .B(_681__31_), .Q(_589_) );
NA2X1 NA2X1_166 ( .gnd!(gnd!), .vdd!(vdd!), .A(_476__bF_buf4), .B(rfRS1[31]), .Q(_590_) );
AN21X1 AN21X1_76 ( .gnd!(gnd!), .vdd!(vdd!), .A(_590_), .B(_473__bF_buf0), .C(_471__bF_buf6), .Q(_591_) );
ON21X1 ON21X1_180 ( .gnd!(gnd!), .vdd!(vdd!), .A(_431_), .B(_473__bF_buf0), .C(_591_), .Q(_592_) );
NA2X1 NA2X1_167 ( .gnd!(gnd!), .vdd!(vdd!), .A(_592_), .B(_589_), .Q(_3__31_) );
MU2X1 MU2X1_80 ( .gnd!(gnd!), .vdd!(vdd!), .IN0(PC1_0_), .IN1(PC_0_), .Q(_2__0_), .S(CTRL_cyc_bF_buf13_bF_buf0) );
MU2X1 MU2X1_81 ( .gnd!(gnd!), .vdd!(vdd!), .IN0(PC1_1_), .IN1(PC_1_), .Q(_2__1_), .S(CTRL_cyc_bF_buf12_bF_buf0) );
MU2X1 MU2X1_82 ( .gnd!(gnd!), .vdd!(vdd!), .IN0(PC1_2_), .IN1(PC_2_), .Q(_2__2_), .S(CTRL_cyc_bF_buf11_bF_buf3) );
MU2X1 MU2X1_83 ( .gnd!(gnd!), .vdd!(vdd!), .IN0(PC1_3_), .IN1(PC_3_), .Q(_2__3_), .S(CTRL_cyc_bF_buf10_bF_buf1) );
MU2X1 MU2X1_84 ( .gnd!(gnd!), .vdd!(vdd!), .IN0(PC1_4_), .IN1(PC_4_), .Q(_2__4_), .S(CTRL_cyc_bF_buf9_bF_buf2) );
MU2IX1 MU2IX1_7 ( .gnd!(gnd!), .vdd!(vdd!), .IN0(_460_), .IN1(_96_), .Q(_2__5_), .S(CTRL_cyc_bF_buf8_bF_buf1) );
MU2X1 MU2X1_85 ( .gnd!(gnd!), .vdd!(vdd!), .IN0(PC1_6_), .IN1(PC_6_), .Q(_2__6_), .S(CTRL_cyc_bF_buf7_bF_buf0) );
MU2X1 MU2X1_86 ( .gnd!(gnd!), .vdd!(vdd!), .IN0(PC1_7_), .IN1(PC_7_), .Q(_2__7_), .S(CTRL_cyc_bF_buf6_bF_buf1) );
MU2IX1 MU2IX1_8 ( .gnd!(gnd!), .vdd!(vdd!), .IN0(_462_), .IN1(_133_), .Q(_2__8_), .S(CTRL_cyc_bF_buf5_bF_buf0) );
MU2X1 MU2X1_87 ( .gnd!(gnd!), .vdd!(vdd!), .IN0(PC1_9_), .IN1(PC_9_), .Q(_2__9_), .S(CTRL_cyc_bF_buf4_bF_buf1) );
MU2X1 MU2X1_88 ( .gnd!(gnd!), .vdd!(vdd!), .IN0(PC1_10_), .IN1(PC_10_), .Q(_2__10_), .S(CTRL_cyc_bF_buf3_bF_buf1) );
MU2X1 MU2X1_89 ( .gnd!(gnd!), .vdd!(vdd!), .IN0(PC1_11_), .IN1(PC_11_), .Q(_2__11_), .S(CTRL_cyc_bF_buf2_bF_buf1) );
MU2X1 MU2X1_90 ( .gnd!(gnd!), .vdd!(vdd!), .IN0(PC1_12_), .IN1(PC_12_), .Q(_2__12_), .S(CTRL_cyc_bF_buf1_bF_buf2) );
MU2X1 MU2X1_91 ( .gnd!(gnd!), .vdd!(vdd!), .IN0(PC1_13_), .IN1(PC_13_), .Q(_2__13_), .S(CTRL_cyc_bF_buf0_bF_buf1) );
MU2X1 MU2X1_92 ( .gnd!(gnd!), .vdd!(vdd!), .IN0(PC1_14_), .IN1(PC_14_), .Q(_2__14_), .S(CTRL_cyc_bF_buf14_bF_buf3) );
MU2X1 MU2X1_93 ( .gnd!(gnd!), .vdd!(vdd!), .IN0(PC1_15_), .IN1(PC_15_), .Q(_2__15_), .S(CTRL_cyc_bF_buf13_bF_buf3) );
MU2IX1 MU2IX1_9 ( .gnd!(gnd!), .vdd!(vdd!), .IN0(_464_), .IN1(_235_), .Q(_2__16_), .S(CTRL_cyc_bF_buf12_bF_buf0) );
MU2X1 MU2X1_94 ( .gnd!(gnd!), .vdd!(vdd!), .IN0(PC1_17_), .IN1(PC_17_), .Q(_2__17_), .S(CTRL_cyc_bF_buf11_bF_buf3) );
MU2X1 MU2X1_95 ( .gnd!(gnd!), .vdd!(vdd!), .IN0(PC1_18_), .IN1(PC_18_), .Q(_2__18_), .S(CTRL_cyc_bF_buf10_bF_buf1) );
MU2X1 MU2X1_96 ( .gnd!(gnd!), .vdd!(vdd!), .IN0(PC1_19_), .IN1(PC_19_), .Q(_2__19_), .S(CTRL_cyc_bF_buf9_bF_buf2) );
MU2IX1 MU2IX1_10 ( .gnd!(gnd!), .vdd!(vdd!), .IN0(_466_), .IN1(_287_), .Q(_2__20_), .S(CTRL_cyc_bF_buf8_bF_buf1) );
MU2IX1 MU2IX1_11 ( .gnd!(gnd!), .vdd!(vdd!), .IN0(_468_), .IN1(_299_), .Q(_2__21_), .S(CTRL_cyc_bF_buf7_bF_buf0) );
MU2X1 MU2X1_97 ( .gnd!(gnd!), .vdd!(vdd!), .IN0(PC1_22_), .IN1(PC_22_), .Q(_2__22_), .S(CTRL_cyc_bF_buf6_bF_buf3) );
MU2X1 MU2X1_98 ( .gnd!(gnd!), .vdd!(vdd!), .IN0(PC1_23_), .IN1(PC_23_), .Q(_2__23_), .S(CTRL_cyc_bF_buf5_bF_buf0) );
MU2X1 MU2X1_99 ( .gnd!(gnd!), .vdd!(vdd!), .IN0(PC1_24_), .IN1(PC_24_), .Q(_2__24_), .S(CTRL_cyc_bF_buf4_bF_buf3) );
MU2X1 MU2X1_100 ( .gnd!(gnd!), .vdd!(vdd!), .IN0(PC1_25_), .IN1(PC_25_), .Q(_2__25_), .S(CTRL_cyc_bF_buf3_bF_buf1) );
MU2X1 MU2X1_101 ( .gnd!(gnd!), .vdd!(vdd!), .IN0(PC1_26_), .IN1(PC_26_), .Q(_2__26_), .S(CTRL_cyc_bF_buf2_bF_buf1) );
MU2X1 MU2X1_102 ( .gnd!(gnd!), .vdd!(vdd!), .IN0(PC1_27_), .IN1(PC_27_), .Q(_2__27_), .S(CTRL_cyc_bF_buf1_bF_buf1) );
MU2IX1 MU2IX1_12 ( .gnd!(gnd!), .vdd!(vdd!), .IN0(_470_), .IN1(_388_), .Q(_2__28_), .S(CTRL_cyc_bF_buf0_bF_buf1) );
MU2X1 MU2X1_103 ( .gnd!(gnd!), .vdd!(vdd!), .IN0(PC1_29_), .IN1(PC_29_), .Q(_2__29_), .S(CTRL_cyc_bF_buf14_bF_buf3) );
MU2X1 MU2X1_104 ( .gnd!(gnd!), .vdd!(vdd!), .IN0(PC1_30_), .IN1(PC_30_), .Q(_2__30_), .S(CTRL_cyc_bF_buf13_bF_buf0) );
MU2X1 MU2X1_105 ( .gnd!(gnd!), .vdd!(vdd!), .IN0(PC1_31_), .IN1(PC_31_), .Q(_2__31_), .S(CTRL_cyc_bF_buf12_bF_buf2) );
MU2X1 MU2X1_106 ( .gnd!(gnd!), .vdd!(vdd!), .IN0(I1_0_), .IN1(IMM_0_), .Q(_0__0_), .S(CTRL_cyc_bF_buf11_bF_buf1) );
MU2X1 MU2X1_107 ( .gnd!(gnd!), .vdd!(vdd!), .IN0(I1_1_), .IN1(IMM_1_), .Q(_0__1_), .S(CTRL_cyc_bF_buf10_bF_buf1) );
MU2X1 MU2X1_108 ( .gnd!(gnd!), .vdd!(vdd!), .IN0(I1_2_), .IN1(IMM_2_), .Q(_0__2_), .S(CTRL_cyc_bF_buf9_bF_buf2) );
MU2X1 MU2X1_109 ( .gnd!(gnd!), .vdd!(vdd!), .IN0(I1_3_), .IN1(IMM_3_), .Q(_0__3_), .S(CTRL_cyc_bF_buf8_bF_buf0) );
MU2X1 MU2X1_110 ( .gnd!(gnd!), .vdd!(vdd!), .IN0(I1_4_), .IN1(IMM_4_), .Q(_0__4_), .S(CTRL_cyc_bF_buf7_bF_buf3) );
MU2X1 MU2X1_111 ( .gnd!(gnd!), .vdd!(vdd!), .IN0(I1_5_), .IN1(IMM_5_), .Q(_0__5_), .S(CTRL_cyc_bF_buf6_bF_buf1) );
MU2X1 MU2X1_112 ( .gnd!(gnd!), .vdd!(vdd!), .IN0(I1_6_), .IN1(IMM_6_), .Q(_0__6_), .S(CTRL_cyc_bF_buf5_bF_buf0) );
MU2X1 MU2X1_113 ( .gnd!(gnd!), .vdd!(vdd!), .IN0(I1_7_), .IN1(IMM_7_), .Q(_0__7_), .S(CTRL_cyc_bF_buf4_bF_buf3) );
MU2X1 MU2X1_114 ( .gnd!(gnd!), .vdd!(vdd!), .IN0(I1_8_), .IN1(IMM_8_), .Q(_0__8_), .S(CTRL_cyc_bF_buf3_bF_buf2) );
MU2X1 MU2X1_115 ( .gnd!(gnd!), .vdd!(vdd!), .IN0(I1_9_), .IN1(IMM_9_), .Q(_0__9_), .S(CTRL_cyc_bF_buf2_bF_buf3) );
MU2X1 MU2X1_116 ( .gnd!(gnd!), .vdd!(vdd!), .IN0(I1_10_), .IN1(IMM_10_), .Q(_0__10_), .S(CTRL_cyc_bF_buf1_bF_buf1) );
MU2X1 MU2X1_117 ( .gnd!(gnd!), .vdd!(vdd!), .IN0(I1_11_), .IN1(IMM_11_), .Q(_0__11_), .S(CTRL_cyc_bF_buf0_bF_buf1) );
MU2X1 MU2X1_118 ( .gnd!(gnd!), .vdd!(vdd!), .IN0(I1_12_), .IN1(IMM_12_), .Q(_0__12_), .S(CTRL_cyc_bF_buf14_bF_buf3) );
MU2X1 MU2X1_119 ( .gnd!(gnd!), .vdd!(vdd!), .IN0(I1_13_), .IN1(IMM_13_), .Q(_0__13_), .S(CTRL_cyc_bF_buf13_bF_buf3) );
MU2X1 MU2X1_120 ( .gnd!(gnd!), .vdd!(vdd!), .IN0(I1_14_), .IN1(IMM_14_), .Q(_0__14_), .S(CTRL_cyc_bF_buf12_bF_buf2) );
MU2X1 MU2X1_121 ( .gnd!(gnd!), .vdd!(vdd!), .IN0(I1_15_), .IN1(IMM_15_), .Q(_0__15_), .S(CTRL_cyc_bF_buf11_bF_buf3) );
MU2X1 MU2X1_122 ( .gnd!(gnd!), .vdd!(vdd!), .IN0(I1_16_), .IN1(IMM_16_), .Q(_0__16_), .S(CTRL_cyc_bF_buf10_bF_buf1) );
MU2X1 MU2X1_123 ( .gnd!(gnd!), .vdd!(vdd!), .IN0(I1_17_), .IN1(IMM_17_), .Q(_0__17_), .S(CTRL_cyc_bF_buf9_bF_buf2) );
MU2X1 MU2X1_124 ( .gnd!(gnd!), .vdd!(vdd!), .IN0(I1_18_), .IN1(IMM_18_), .Q(_0__18_), .S(CTRL_cyc_bF_buf8_bF_buf0) );
MU2X1 MU2X1_125 ( .gnd!(gnd!), .vdd!(vdd!), .IN0(I1_19_), .IN1(IMM_19_), .Q(_0__19_), .S(CTRL_cyc_bF_buf7_bF_buf2) );
MU2X1 MU2X1_126 ( .gnd!(gnd!), .vdd!(vdd!), .IN0(I1_20_), .IN1(IMM_20_), .Q(_0__20_), .S(CTRL_cyc_bF_buf6_bF_buf3) );
MU2X1 MU2X1_127 ( .gnd!(gnd!), .vdd!(vdd!), .IN0(I1_21_), .IN1(IMM_21_), .Q(_0__21_), .S(CTRL_cyc_bF_buf5_bF_buf1) );
MU2X1 MU2X1_128 ( .gnd!(gnd!), .vdd!(vdd!), .IN0(I1_22_), .IN1(IMM_22_), .Q(_0__22_), .S(CTRL_cyc_bF_buf4_bF_buf3) );
MU2X1 MU2X1_129 ( .gnd!(gnd!), .vdd!(vdd!), .IN0(I1_23_), .IN1(IMM_23_), .Q(_0__23_), .S(CTRL_cyc_bF_buf3_bF_buf1) );
MU2X1 MU2X1_130 ( .gnd!(gnd!), .vdd!(vdd!), .IN0(I1_24_), .IN1(IMM_24_), .Q(_0__24_), .S(CTRL_cyc_bF_buf2_bF_buf3) );
MU2X1 MU2X1_131 ( .gnd!(gnd!), .vdd!(vdd!), .IN0(I1_25_), .IN1(IMM_25_), .Q(_0__25_), .S(CTRL_cyc_bF_buf1_bF_buf1) );
MU2X1 MU2X1_132 ( .gnd!(gnd!), .vdd!(vdd!), .IN0(I1_26_), .IN1(IMM_26_), .Q(_0__26_), .S(CTRL_cyc_bF_buf0_bF_buf1) );
MU2X1 MU2X1_133 ( .gnd!(gnd!), .vdd!(vdd!), .IN0(I1_27_), .IN1(IMM_27_), .Q(_0__27_), .S(CTRL_cyc_bF_buf14_bF_buf2) );
MU2X1 MU2X1_134 ( .gnd!(gnd!), .vdd!(vdd!), .IN0(I1_28_), .IN1(IMM_28_), .Q(_0__28_), .S(CTRL_cyc_bF_buf13_bF_buf2) );
MU2X1 MU2X1_135 ( .gnd!(gnd!), .vdd!(vdd!), .IN0(I1_29_), .IN1(IMM_29_), .Q(_0__29_), .S(CTRL_cyc_bF_buf12_bF_buf2) );
MU2X1 MU2X1_136 ( .gnd!(gnd!), .vdd!(vdd!), .IN0(I1_30_), .IN1(IMM_30_), .Q(_0__30_), .S(CTRL_cyc_bF_buf11_bF_buf3) );
MU2X1 MU2X1_137 ( .gnd!(gnd!), .vdd!(vdd!), .IN0(I1_31_), .IN1(CTRL_IDEC0_IR_31_), .Q(_0__31_), .S(CTRL_cyc_bF_buf10_bF_buf0) );
MU2X1 MU2X1_138 ( .gnd!(gnd!), .vdd!(vdd!), .IN0(bdo[0]), .IN1(CTRL_IDEC0_IR_0_), .Q(_1__0_), .S(CTRL_cyc_bF_buf9_bF_buf1) );
MU2X1 MU2X1_139 ( .gnd!(gnd!), .vdd!(vdd!), .IN0(bdo[1]), .IN1(CTRL_IDEC0_IR_1_), .Q(_1__1_), .S(CTRL_cyc_bF_buf8_bF_buf2) );
MU2X1 MU2X1_140 ( .gnd!(gnd!), .vdd!(vdd!), .IN0(bdo[2]), .IN1(CTRL_IDEC0_IR_2_), .Q(_1__2_), .S(CTRL_cyc_bF_buf7_bF_buf3) );
MU2X1 MU2X1_141 ( .gnd!(gnd!), .vdd!(vdd!), .IN0(bdo[3]), .IN1(CTRL_IDEC0_IR_3_), .Q(_1__3_), .S(CTRL_cyc_bF_buf6_bF_buf2) );
MU2X1 MU2X1_142 ( .gnd!(gnd!), .vdd!(vdd!), .IN0(bdo[4]), .IN1(CTRL_IDEC0_IR_4_), .Q(_1__4_), .S(CTRL_cyc_bF_buf5_bF_buf3) );
MU2X1 MU2X1_143 ( .gnd!(gnd!), .vdd!(vdd!), .IN0(bdo[5]), .IN1(CTRL_IDEC0_IR_5_), .Q(_1__5_), .S(CTRL_cyc_bF_buf4_bF_buf1) );
MU2X1 MU2X1_144 ( .gnd!(gnd!), .vdd!(vdd!), .IN0(bdo[6]), .IN1(CTRL_IDEC0_IR_6_), .Q(_1__6_), .S(CTRL_cyc_bF_buf3_bF_buf2) );
MU2X1 MU2X1_145 ( .gnd!(gnd!), .vdd!(vdd!), .IN0(bdo[7]), .IN1(CTRL_IDEC0_IR_7_), .Q(_1__7_), .S(CTRL_cyc_bF_buf2_bF_buf0) );
MU2X1 MU2X1_146 ( .gnd!(gnd!), .vdd!(vdd!), .IN0(bdo[8]), .IN1(CTRL_IDEC0_IR_8_), .Q(_1__8_), .S(CTRL_cyc_bF_buf1_bF_buf1) );
MU2X1 MU2X1_147 ( .gnd!(gnd!), .vdd!(vdd!), .IN0(bdo[9]), .IN1(CTRL_IDEC0_IR_9_), .Q(_1__9_), .S(CTRL_cyc_bF_buf0_bF_buf3) );
MU2X1 MU2X1_148 ( .gnd!(gnd!), .vdd!(vdd!), .IN0(bdo[10]), .IN1(CTRL_IDEC0_IR_10_), .Q(_1__10_), .S(CTRL_cyc_bF_buf14_bF_buf2) );
MU2X1 MU2X1_149 ( .gnd!(gnd!), .vdd!(vdd!), .IN0(bdo[11]), .IN1(CTRL_IDEC0_IR_11_), .Q(_1__11_), .S(CTRL_cyc_bF_buf13_bF_buf3) );
MU2X1 MU2X1_150 ( .gnd!(gnd!), .vdd!(vdd!), .IN0(bdo[12]), .IN1(CTRL_IDEC0_IR_12_), .Q(_1__12_), .S(CTRL_cyc_bF_buf12_bF_buf3) );
MU2X1 MU2X1_151 ( .gnd!(gnd!), .vdd!(vdd!), .IN0(bdo[13]), .IN1(CTRL_IDEC0_IR_13_), .Q(_1__13_), .S(CTRL_cyc_bF_buf11_bF_buf2) );
MU2X1 MU2X1_152 ( .gnd!(gnd!), .vdd!(vdd!), .IN0(bdo[14]), .IN1(CTRL_IDEC0_IR_14_), .Q(_1__14_), .S(CTRL_cyc_bF_buf10_bF_buf3) );
MU2X1 MU2X1_153 ( .gnd!(gnd!), .vdd!(vdd!), .IN0(bdo[15]), .IN1(_686__0_), .Q(_1__15_), .S(CTRL_cyc_bF_buf9_bF_buf3) );
MU2X1 MU2X1_154 ( .gnd!(gnd!), .vdd!(vdd!), .IN0(bdo[16]), .IN1(_686__1_), .Q(_1__16_), .S(CTRL_cyc_bF_buf8_bF_buf3) );
MU2X1 MU2X1_155 ( .gnd!(gnd!), .vdd!(vdd!), .IN0(bdo[17]), .IN1(_686__2_), .Q(_1__17_), .S(CTRL_cyc_bF_buf7_bF_buf1) );
MU2X1 MU2X1_156 ( .gnd!(gnd!), .vdd!(vdd!), .IN0(bdo[18]), .IN1(_686__3_), .Q(_1__18_), .S(CTRL_cyc_bF_buf6_bF_buf2) );
MU2X1 MU2X1_157 ( .gnd!(gnd!), .vdd!(vdd!), .IN0(bdo[19]), .IN1(_686__4_), .Q(_1__19_), .S(CTRL_cyc_bF_buf5_bF_buf3) );
MU2X1 MU2X1_158 ( .gnd!(gnd!), .vdd!(vdd!), .IN0(bdo[20]), .IN1(_687__0_), .Q(_1__20_), .S(CTRL_cyc_bF_buf4_bF_buf2) );
MU2X1 MU2X1_159 ( .gnd!(gnd!), .vdd!(vdd!), .IN0(bdo[21]), .IN1(_687__1_), .Q(_1__21_), .S(CTRL_cyc_bF_buf3_bF_buf0) );
MU2X1 MU2X1_160 ( .gnd!(gnd!), .vdd!(vdd!), .IN0(bdo[22]), .IN1(_687__2_), .Q(_1__22_), .S(CTRL_cyc_bF_buf2_bF_buf0) );
MU2X1 MU2X1_161 ( .gnd!(gnd!), .vdd!(vdd!), .IN0(bdo[23]), .IN1(_687__3_), .Q(_1__23_), .S(CTRL_cyc_bF_buf1_bF_buf3) );
MU2X1 MU2X1_162 ( .gnd!(gnd!), .vdd!(vdd!), .IN0(bdo[24]), .IN1(_687__4_), .Q(_1__24_), .S(CTRL_cyc_bF_buf0_bF_buf3) );
MU2X1 MU2X1_163 ( .gnd!(gnd!), .vdd!(vdd!), .IN0(bdo[25]), .IN1(CTRL_IDEC0_IR_25_), .Q(_1__25_), .S(CTRL_cyc_bF_buf14_bF_buf1) );
MU2X1 MU2X1_164 ( .gnd!(gnd!), .vdd!(vdd!), .IN0(bdo[26]), .IN1(CTRL_IDEC0_IR_26_), .Q(_1__26_), .S(CTRL_cyc_bF_buf13_bF_buf2) );
MU2X1 MU2X1_165 ( .gnd!(gnd!), .vdd!(vdd!), .IN0(bdo[27]), .IN1(CTRL_IDEC0_IR_27_), .Q(_1__27_), .S(CTRL_cyc_bF_buf12_bF_buf3) );
MU2X1 MU2X1_166 ( .gnd!(gnd!), .vdd!(vdd!), .IN0(bdo[28]), .IN1(CTRL_IDEC0_IR_28_), .Q(_1__28_), .S(CTRL_cyc_bF_buf11_bF_buf2) );
MU2X1 MU2X1_167 ( .gnd!(gnd!), .vdd!(vdd!), .IN0(bdo[29]), .IN1(CTRL_IDEC0_IR_29_), .Q(_1__29_), .S(CTRL_cyc_bF_buf10_bF_buf0) );
MU2X1 MU2X1_168 ( .gnd!(gnd!), .vdd!(vdd!), .IN0(bdo[30]), .IN1(CTRL_IDEC0_IR_30_), .Q(_1__30_), .S(CTRL_cyc_bF_buf9_bF_buf3) );
MU2X1 MU2X1_169 ( .gnd!(gnd!), .vdd!(vdd!), .IN0(bdo[31]), .IN1(CTRL_IDEC0_IR_31_), .Q(_1__31_), .S(CTRL_cyc_bF_buf8_bF_buf3) );
INX4 INX4_1 ( .gnd!(gnd!), .vdd!(vdd!), .A(rst), .Q(_268_) );
BUX1 BUX1_1 ( .gnd!(gnd!), .vdd!(vdd!), .A(_677__0_), .Q(baddr[0]) );
BUX1 BUX1_2 ( .gnd!(gnd!), .vdd!(vdd!), .A(_677__1_), .Q(baddr[1]) );
BUX1 BUX1_3 ( .gnd!(gnd!), .vdd!(vdd!), .A(_677__2_), .Q(baddr[2]) );
BUX1 BUX1_4 ( .gnd!(gnd!), .vdd!(vdd!), .A(_677__3_), .Q(baddr[3]) );
BUX1 BUX1_5 ( .gnd!(gnd!), .vdd!(vdd!), .A(_677__4_), .Q(baddr[4]) );
BUX1 BUX1_6 ( .gnd!(gnd!), .vdd!(vdd!), .A(_677__5_), .Q(baddr[5]) );
BUX1 BUX1_7 ( .gnd!(gnd!), .vdd!(vdd!), .A(_677__6_), .Q(baddr[6]) );
BUX1 BUX1_8 ( .gnd!(gnd!), .vdd!(vdd!), .A(_677__7_), .Q(baddr[7]) );
BUX1 BUX1_9 ( .gnd!(gnd!), .vdd!(vdd!), .A(_677__8_), .Q(baddr[8]) );
BUX1 BUX1_10 ( .gnd!(gnd!), .vdd!(vdd!), .A(_677__9_), .Q(baddr[9]) );
BUX1 BUX1_11 ( .gnd!(gnd!), .vdd!(vdd!), .A(_677__10_), .Q(baddr[10]) );
BUX1 BUX1_12 ( .gnd!(gnd!), .vdd!(vdd!), .A(_677__11_), .Q(baddr[11]) );
BUX1 BUX1_13 ( .gnd!(gnd!), .vdd!(vdd!), .A(_677__12_), .Q(baddr[12]) );
BUX1 BUX1_14 ( .gnd!(gnd!), .vdd!(vdd!), .A(_677__13_), .Q(baddr[13]) );
BUX1 BUX1_15 ( .gnd!(gnd!), .vdd!(vdd!), .A(_677__14_), .Q(baddr[14]) );
BUX1 BUX1_16 ( .gnd!(gnd!), .vdd!(vdd!), .A(_677__15_), .Q(baddr[15]) );
BUX1 BUX1_17 ( .gnd!(gnd!), .vdd!(vdd!), .A(_677__16_), .Q(baddr[16]) );
BUX1 BUX1_18 ( .gnd!(gnd!), .vdd!(vdd!), .A(_677__17_), .Q(baddr[17]) );
BUX1 BUX1_19 ( .gnd!(gnd!), .vdd!(vdd!), .A(_677__18_), .Q(baddr[18]) );
BUX1 BUX1_20 ( .gnd!(gnd!), .vdd!(vdd!), .A(_677__19_), .Q(baddr[19]) );
BUX1 BUX1_21 ( .gnd!(gnd!), .vdd!(vdd!), .A(_677__20_), .Q(baddr[20]) );
BUX1 BUX1_22 ( .gnd!(gnd!), .vdd!(vdd!), .A(_677__21_), .Q(baddr[21]) );
BUX1 BUX1_23 ( .gnd!(gnd!), .vdd!(vdd!), .A(_677__22_), .Q(baddr[22]) );
BUX1 BUX1_24 ( .gnd!(gnd!), .vdd!(vdd!), .A(_677__23_), .Q(baddr[23]) );
BUX1 BUX1_25 ( .gnd!(gnd!), .vdd!(vdd!), .A(_677__24_), .Q(baddr[24]) );
BUX1 BUX1_26 ( .gnd!(gnd!), .vdd!(vdd!), .A(_677__25_), .Q(baddr[25]) );
BUX1 BUX1_27 ( .gnd!(gnd!), .vdd!(vdd!), .A(_677__26_), .Q(baddr[26]) );
BUX1 BUX1_28 ( .gnd!(gnd!), .vdd!(vdd!), .A(_677__27_), .Q(baddr[27]) );
BUX1 BUX1_29 ( .gnd!(gnd!), .vdd!(vdd!), .A(_677__28_), .Q(baddr[28]) );
BUX1 BUX1_30 ( .gnd!(gnd!), .vdd!(vdd!), .A(_677__29_), .Q(baddr[29]) );
BUX1 BUX1_31 ( .gnd!(gnd!), .vdd!(vdd!), .A(_677__30_), .Q(baddr[30]) );
BUX1 BUX1_32 ( .gnd!(gnd!), .vdd!(vdd!), .A(_677__31_), .Q(baddr[31]) );
BUX1 BUX1_33 ( .gnd!(gnd!), .vdd!(vdd!), .A(_678__0_), .Q(bdi[0]) );
BUX1 BUX1_34 ( .gnd!(gnd!), .vdd!(vdd!), .A(_678__1_), .Q(bdi[1]) );
BUX1 BUX1_35 ( .gnd!(gnd!), .vdd!(vdd!), .A(_678__2_), .Q(bdi[2]) );
BUX1 BUX1_36 ( .gnd!(gnd!), .vdd!(vdd!), .A(_678__3_), .Q(bdi[3]) );
BUX1 BUX1_37 ( .gnd!(gnd!), .vdd!(vdd!), .A(_678__4_), .Q(bdi[4]) );
BUX1 BUX1_38 ( .gnd!(gnd!), .vdd!(vdd!), .A(_678__5_), .Q(bdi[5]) );
BUX1 BUX1_39 ( .gnd!(gnd!), .vdd!(vdd!), .A(_678__6_), .Q(bdi[6]) );
BUX1 BUX1_40 ( .gnd!(gnd!), .vdd!(vdd!), .A(_678__7_), .Q(bdi[7]) );
BUX1 BUX1_41 ( .gnd!(gnd!), .vdd!(vdd!), .A(_678__8_), .Q(bdi[8]) );
BUX1 BUX1_42 ( .gnd!(gnd!), .vdd!(vdd!), .A(_678__9_), .Q(bdi[9]) );
BUX1 BUX1_43 ( .gnd!(gnd!), .vdd!(vdd!), .A(_678__10_), .Q(bdi[10]) );
BUX1 BUX1_44 ( .gnd!(gnd!), .vdd!(vdd!), .A(_678__11_), .Q(bdi[11]) );
BUX1 BUX1_45 ( .gnd!(gnd!), .vdd!(vdd!), .A(_678__12_), .Q(bdi[12]) );
BUX1 BUX1_46 ( .gnd!(gnd!), .vdd!(vdd!), .A(_678__13_), .Q(bdi[13]) );
BUX1 BUX1_47 ( .gnd!(gnd!), .vdd!(vdd!), .A(_678__14_), .Q(bdi[14]) );
BUX1 BUX1_48 ( .gnd!(gnd!), .vdd!(vdd!), .A(_678__15_), .Q(bdi[15]) );
BUX1 BUX1_49 ( .gnd!(gnd!), .vdd!(vdd!), .A(_678__16_), .Q(bdi[16]) );
BUX1 BUX1_50 ( .gnd!(gnd!), .vdd!(vdd!), .A(_678__17_), .Q(bdi[17]) );
BUX1 BUX1_51 ( .gnd!(gnd!), .vdd!(vdd!), .A(_678__18_), .Q(bdi[18]) );
BUX1 BUX1_52 ( .gnd!(gnd!), .vdd!(vdd!), .A(_678__19_), .Q(bdi[19]) );
BUX1 BUX1_53 ( .gnd!(gnd!), .vdd!(vdd!), .A(_678__20_), .Q(bdi[20]) );
BUX1 BUX1_54 ( .gnd!(gnd!), .vdd!(vdd!), .A(_678__21_), .Q(bdi[21]) );
BUX1 BUX1_55 ( .gnd!(gnd!), .vdd!(vdd!), .A(_678__22_), .Q(bdi[22]) );
BUX1 BUX1_56 ( .gnd!(gnd!), .vdd!(vdd!), .A(_678__23_), .Q(bdi[23]) );
BUX1 BUX1_57 ( .gnd!(gnd!), .vdd!(vdd!), .A(_678__24_), .Q(bdi[24]) );
BUX1 BUX1_58 ( .gnd!(gnd!), .vdd!(vdd!), .A(_678__25_), .Q(bdi[25]) );
BUX1 BUX1_59 ( .gnd!(gnd!), .vdd!(vdd!), .A(_678__26_), .Q(bdi[26]) );
BUX1 BUX1_60 ( .gnd!(gnd!), .vdd!(vdd!), .A(_678__27_), .Q(bdi[27]) );
BUX1 BUX1_61 ( .gnd!(gnd!), .vdd!(vdd!), .A(_678__28_), .Q(bdi[28]) );
BUX1 BUX1_62 ( .gnd!(gnd!), .vdd!(vdd!), .A(_678__29_), .Q(bdi[29]) );
BUX1 BUX1_63 ( .gnd!(gnd!), .vdd!(vdd!), .A(_678__30_), .Q(bdi[30]) );
BUX1 BUX1_64 ( .gnd!(gnd!), .vdd!(vdd!), .A(_678__31_), .Q(bdi[31]) );
BUX1 BUX1_65 ( .gnd!(gnd!), .vdd!(vdd!), .A(_679__0_), .Q(bsz[0]) );
BUX1 BUX1_66 ( .gnd!(gnd!), .vdd!(vdd!), .A(_679__1_), .Q(bsz[1]) );
BUX1 BUX1_67 ( .gnd!(gnd!), .vdd!(vdd!), .A(_680_), .Q(bwr) );
BUX1 BUX1_68 ( .gnd!(gnd!), .vdd!(vdd!), .A(_681__0_), .Q(extA[0]) );
BUX1 BUX1_69 ( .gnd!(gnd!), .vdd!(vdd!), .A(_681__1_), .Q(extA[1]) );
BUX1 BUX1_70 ( .gnd!(gnd!), .vdd!(vdd!), .A(_681__2_), .Q(extA[2]) );
BUX1 BUX1_71 ( .gnd!(gnd!), .vdd!(vdd!), .A(_681__3_), .Q(extA[3]) );
BUX1 BUX1_72 ( .gnd!(gnd!), .vdd!(vdd!), .A(_681__4_), .Q(extA[4]) );
BUX1 BUX1_73 ( .gnd!(gnd!), .vdd!(vdd!), .A(_681__5_), .Q(extA[5]) );
BUX1 BUX1_74 ( .gnd!(gnd!), .vdd!(vdd!), .A(_681__6_), .Q(extA[6]) );
BUX1 BUX1_75 ( .gnd!(gnd!), .vdd!(vdd!), .A(_681__7_), .Q(extA[7]) );
BUX1 BUX1_76 ( .gnd!(gnd!), .vdd!(vdd!), .A(_681__8_), .Q(extA[8]) );
BUX1 BUX1_77 ( .gnd!(gnd!), .vdd!(vdd!), .A(_681__9_), .Q(extA[9]) );
BUX1 BUX1_78 ( .gnd!(gnd!), .vdd!(vdd!), .A(_681__10_), .Q(extA[10]) );
BUX1 BUX1_79 ( .gnd!(gnd!), .vdd!(vdd!), .A(_681__11_), .Q(extA[11]) );
BUX1 BUX1_80 ( .gnd!(gnd!), .vdd!(vdd!), .A(_681__12_), .Q(extA[12]) );
BUX1 BUX1_81 ( .gnd!(gnd!), .vdd!(vdd!), .A(_681__13_), .Q(extA[13]) );
BUX1 BUX1_82 ( .gnd!(gnd!), .vdd!(vdd!), .A(_681__14_), .Q(extA[14]) );
BUX1 BUX1_83 ( .gnd!(gnd!), .vdd!(vdd!), .A(_681__15_), .Q(extA[15]) );
BUX1 BUX1_84 ( .gnd!(gnd!), .vdd!(vdd!), .A(_681__16_), .Q(extA[16]) );
BUX1 BUX1_85 ( .gnd!(gnd!), .vdd!(vdd!), .A(_681__17_), .Q(extA[17]) );
BUX1 BUX1_86 ( .gnd!(gnd!), .vdd!(vdd!), .A(_681__18_), .Q(extA[18]) );
BUX1 BUX1_87 ( .gnd!(gnd!), .vdd!(vdd!), .A(_681__19_), .Q(extA[19]) );
BUX1 BUX1_88 ( .gnd!(gnd!), .vdd!(vdd!), .A(_681__20_), .Q(extA[20]) );
BUX1 BUX1_89 ( .gnd!(gnd!), .vdd!(vdd!), .A(_681__21_), .Q(extA[21]) );
BUX1 BUX1_90 ( .gnd!(gnd!), .vdd!(vdd!), .A(_681__22_), .Q(extA[22]) );
BUX1 BUX1_91 ( .gnd!(gnd!), .vdd!(vdd!), .A(_681__23_), .Q(extA[23]) );
BUX1 BUX1_92 ( .gnd!(gnd!), .vdd!(vdd!), .A(_681__24_), .Q(extA[24]) );
BUX1 BUX1_93 ( .gnd!(gnd!), .vdd!(vdd!), .A(_681__25_), .Q(extA[25]) );
BUX1 BUX1_94 ( .gnd!(gnd!), .vdd!(vdd!), .A(_681__26_), .Q(extA[26]) );
BUX1 BUX1_95 ( .gnd!(gnd!), .vdd!(vdd!), .A(_681__27_), .Q(extA[27]) );
BUX1 BUX1_96 ( .gnd!(gnd!), .vdd!(vdd!), .A(_681__28_), .Q(extA[28]) );
BUX1 BUX1_97 ( .gnd!(gnd!), .vdd!(vdd!), .A(_681__29_), .Q(extA[29]) );
BUX1 BUX1_98 ( .gnd!(gnd!), .vdd!(vdd!), .A(_681__30_), .Q(extA[30]) );
BUX1 BUX1_99 ( .gnd!(gnd!), .vdd!(vdd!), .A(_681__31_), .Q(extA[31]) );
BUX1 BUX1_100 ( .gnd!(gnd!), .vdd!(vdd!), .A(_678__0_), .Q(extB[0]) );
BUX1 BUX1_101 ( .gnd!(gnd!), .vdd!(vdd!), .A(_678__1_), .Q(extB[1]) );
BUX1 BUX1_102 ( .gnd!(gnd!), .vdd!(vdd!), .A(_678__2_), .Q(extB[2]) );
BUX1 BUX1_103 ( .gnd!(gnd!), .vdd!(vdd!), .A(_678__3_), .Q(extB[3]) );
BUX1 BUX1_104 ( .gnd!(gnd!), .vdd!(vdd!), .A(_678__4_), .Q(extB[4]) );
BUX1 BUX1_105 ( .gnd!(gnd!), .vdd!(vdd!), .A(_678__5_), .Q(extB[5]) );
BUX1 BUX1_106 ( .gnd!(gnd!), .vdd!(vdd!), .A(_678__6_), .Q(extB[6]) );
BUX1 BUX1_107 ( .gnd!(gnd!), .vdd!(vdd!), .A(_678__7_), .Q(extB[7]) );
BUX1 BUX1_108 ( .gnd!(gnd!), .vdd!(vdd!), .A(_678__8_), .Q(extB[8]) );
BUX1 BUX1_109 ( .gnd!(gnd!), .vdd!(vdd!), .A(_678__9_), .Q(extB[9]) );
BUX1 BUX1_110 ( .gnd!(gnd!), .vdd!(vdd!), .A(_678__10_), .Q(extB[10]) );
BUX1 BUX1_111 ( .gnd!(gnd!), .vdd!(vdd!), .A(_678__11_), .Q(extB[11]) );
BUX1 BUX1_112 ( .gnd!(gnd!), .vdd!(vdd!), .A(_678__12_), .Q(extB[12]) );
BUX1 BUX1_113 ( .gnd!(gnd!), .vdd!(vdd!), .A(_678__13_), .Q(extB[13]) );
BUX1 BUX1_114 ( .gnd!(gnd!), .vdd!(vdd!), .A(_678__14_), .Q(extB[14]) );
BUX1 BUX1_115 ( .gnd!(gnd!), .vdd!(vdd!), .A(_678__15_), .Q(extB[15]) );
BUX1 BUX1_116 ( .gnd!(gnd!), .vdd!(vdd!), .A(_678__16_), .Q(extB[16]) );
BUX1 BUX1_117 ( .gnd!(gnd!), .vdd!(vdd!), .A(_678__17_), .Q(extB[17]) );
BUX1 BUX1_118 ( .gnd!(gnd!), .vdd!(vdd!), .A(_678__18_), .Q(extB[18]) );
BUX1 BUX1_119 ( .gnd!(gnd!), .vdd!(vdd!), .A(_678__19_), .Q(extB[19]) );
BUX1 BUX1_120 ( .gnd!(gnd!), .vdd!(vdd!), .A(_678__20_), .Q(extB[20]) );
BUX1 BUX1_121 ( .gnd!(gnd!), .vdd!(vdd!), .A(_678__21_), .Q(extB[21]) );
BUX1 BUX1_122 ( .gnd!(gnd!), .vdd!(vdd!), .A(_678__22_), .Q(extB[22]) );
BUX1 BUX1_123 ( .gnd!(gnd!), .vdd!(vdd!), .A(_678__23_), .Q(extB[23]) );
BUX1 BUX1_124 ( .gnd!(gnd!), .vdd!(vdd!), .A(_678__24_), .Q(extB[24]) );
BUX1 BUX1_125 ( .gnd!(gnd!), .vdd!(vdd!), .A(_678__25_), .Q(extB[25]) );
BUX1 BUX1_126 ( .gnd!(gnd!), .vdd!(vdd!), .A(_678__26_), .Q(extB[26]) );
BUX1 BUX1_127 ( .gnd!(gnd!), .vdd!(vdd!), .A(_678__27_), .Q(extB[27]) );
BUX1 BUX1_128 ( .gnd!(gnd!), .vdd!(vdd!), .A(_678__28_), .Q(extB[28]) );
BUX1 BUX1_129 ( .gnd!(gnd!), .vdd!(vdd!), .A(_678__29_), .Q(extB[29]) );
BUX1 BUX1_130 ( .gnd!(gnd!), .vdd!(vdd!), .A(_678__30_), .Q(extB[30]) );
BUX1 BUX1_131 ( .gnd!(gnd!), .vdd!(vdd!), .A(_678__31_), .Q(extB[31]) );
BUX1 BUX1_132 ( .gnd!(gnd!), .vdd!(vdd!), .A(_682__0_bF_buf3), .Q(extFunc3[0]) );
BUX1 BUX1_133 ( .gnd!(gnd!), .vdd!(vdd!), .A(_682__1_bF_buf4), .Q(extFunc3[1]) );
BUX1 BUX1_134 ( .gnd!(gnd!), .vdd!(vdd!), .A(EXT_type_bF_buf4), .Q(extFunc3[2]) );
BUX1 BUX1_135 ( .gnd!(gnd!), .vdd!(vdd!), .A(_683_), .Q(extStart) );
BUX1 BUX1_136 ( .gnd!(gnd!), .vdd!(vdd!), .A(_684__0_), .Q(rfD[0]) );
BUX1 BUX1_137 ( .gnd!(gnd!), .vdd!(vdd!), .A(_684__1_), .Q(rfD[1]) );
BUX1 BUX1_138 ( .gnd!(gnd!), .vdd!(vdd!), .A(_684__2_), .Q(rfD[2]) );
BUX1 BUX1_139 ( .gnd!(gnd!), .vdd!(vdd!), .A(_684__3_), .Q(rfD[3]) );
BUX1 BUX1_140 ( .gnd!(gnd!), .vdd!(vdd!), .A(_684__4_), .Q(rfD[4]) );
BUX1 BUX1_141 ( .gnd!(gnd!), .vdd!(vdd!), .A(_684__5_), .Q(rfD[5]) );
BUX1 BUX1_142 ( .gnd!(gnd!), .vdd!(vdd!), .A(_684__6_), .Q(rfD[6]) );
BUX1 BUX1_143 ( .gnd!(gnd!), .vdd!(vdd!), .A(_684__7_), .Q(rfD[7]) );
BUX1 BUX1_144 ( .gnd!(gnd!), .vdd!(vdd!), .A(_684__8_), .Q(rfD[8]) );
BUX1 BUX1_145 ( .gnd!(gnd!), .vdd!(vdd!), .A(_684__9_), .Q(rfD[9]) );
BUX1 BUX1_146 ( .gnd!(gnd!), .vdd!(vdd!), .A(_684__10_), .Q(rfD[10]) );
BUX1 BUX1_147 ( .gnd!(gnd!), .vdd!(vdd!), .A(_684__11_), .Q(rfD[11]) );
BUX1 BUX1_148 ( .gnd!(gnd!), .vdd!(vdd!), .A(_684__12_), .Q(rfD[12]) );
BUX1 BUX1_149 ( .gnd!(gnd!), .vdd!(vdd!), .A(_684__13_), .Q(rfD[13]) );
BUX1 BUX1_150 ( .gnd!(gnd!), .vdd!(vdd!), .A(_684__14_), .Q(rfD[14]) );
BUX1 BUX1_151 ( .gnd!(gnd!), .vdd!(vdd!), .A(_684__15_), .Q(rfD[15]) );
BUX1 BUX1_152 ( .gnd!(gnd!), .vdd!(vdd!), .A(_684__16_), .Q(rfD[16]) );
BUX1 BUX1_153 ( .gnd!(gnd!), .vdd!(vdd!), .A(_684__17_), .Q(rfD[17]) );
BUX1 BUX1_154 ( .gnd!(gnd!), .vdd!(vdd!), .A(_684__18_), .Q(rfD[18]) );
BUX1 BUX1_155 ( .gnd!(gnd!), .vdd!(vdd!), .A(_684__19_), .Q(rfD[19]) );
BUX1 BUX1_156 ( .gnd!(gnd!), .vdd!(vdd!), .A(_684__20_), .Q(rfD[20]) );
BUX1 BUX1_157 ( .gnd!(gnd!), .vdd!(vdd!), .A(_684__21_), .Q(rfD[21]) );
BUX1 BUX1_158 ( .gnd!(gnd!), .vdd!(vdd!), .A(_684__22_), .Q(rfD[22]) );
BUX1 BUX1_159 ( .gnd!(gnd!), .vdd!(vdd!), .A(_684__23_), .Q(rfD[23]) );
BUX1 BUX1_160 ( .gnd!(gnd!), .vdd!(vdd!), .A(_684__24_), .Q(rfD[24]) );
BUX1 BUX1_161 ( .gnd!(gnd!), .vdd!(vdd!), .A(_684__25_), .Q(rfD[25]) );
BUX1 BUX1_162 ( .gnd!(gnd!), .vdd!(vdd!), .A(_684__26_), .Q(rfD[26]) );
BUX1 BUX1_163 ( .gnd!(gnd!), .vdd!(vdd!), .A(_684__27_), .Q(rfD[27]) );
BUX1 BUX1_164 ( .gnd!(gnd!), .vdd!(vdd!), .A(_684__28_), .Q(rfD[28]) );
BUX1 BUX1_165 ( .gnd!(gnd!), .vdd!(vdd!), .A(_684__29_), .Q(rfD[29]) );
BUX1 BUX1_166 ( .gnd!(gnd!), .vdd!(vdd!), .A(_684__30_), .Q(rfD[30]) );
BUX1 BUX1_167 ( .gnd!(gnd!), .vdd!(vdd!), .A(_684__31_), .Q(rfD[31]) );
BUX1 BUX1_168 ( .gnd!(gnd!), .vdd!(vdd!), .A(_685__0_), .Q(rfrd[0]) );
BUX1 BUX1_169 ( .gnd!(gnd!), .vdd!(vdd!), .A(_685__1_), .Q(rfrd[1]) );
BUX1 BUX1_170 ( .gnd!(gnd!), .vdd!(vdd!), .A(_685__2_), .Q(rfrd[2]) );
BUX1 BUX1_171 ( .gnd!(gnd!), .vdd!(vdd!), .A(_685__3_), .Q(rfrd[3]) );
BUX1 BUX1_172 ( .gnd!(gnd!), .vdd!(vdd!), .A(_685__4_), .Q(rfrd[4]) );
BUX1 BUX1_173 ( .gnd!(gnd!), .vdd!(vdd!), .A(_686__0_), .Q(rfrs1[0]) );
BUX1 BUX1_174 ( .gnd!(gnd!), .vdd!(vdd!), .A(_686__1_), .Q(rfrs1[1]) );
BUX1 BUX1_175 ( .gnd!(gnd!), .vdd!(vdd!), .A(_686__2_), .Q(rfrs1[2]) );
BUX1 BUX1_176 ( .gnd!(gnd!), .vdd!(vdd!), .A(_686__3_), .Q(rfrs1[3]) );
BUX1 BUX1_177 ( .gnd!(gnd!), .vdd!(vdd!), .A(_686__4_), .Q(rfrs1[4]) );
BUX1 BUX1_178 ( .gnd!(gnd!), .vdd!(vdd!), .A(_687__0_), .Q(rfrs2[0]) );
BUX1 BUX1_179 ( .gnd!(gnd!), .vdd!(vdd!), .A(_687__1_), .Q(rfrs2[1]) );
BUX1 BUX1_180 ( .gnd!(gnd!), .vdd!(vdd!), .A(_687__2_), .Q(rfrs2[2]) );
BUX1 BUX1_181 ( .gnd!(gnd!), .vdd!(vdd!), .A(_687__3_), .Q(rfrs2[3]) );
BUX1 BUX1_182 ( .gnd!(gnd!), .vdd!(vdd!), .A(_687__4_), .Q(rfrs2[4]) );
BUX1 BUX1_183 ( .gnd!(gnd!), .vdd!(vdd!), .A(_688_), .Q(rfwr) );
DFRQX1 DFRQX1_1 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf14), .D(_6__0_), .Q(R_0_) );
DFRQX1 DFRQX1_2 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf21), .D(_6__1_), .Q(R_1_) );
DFRQX1 DFRQX1_3 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf53), .D(_6__2_), .Q(R_2_) );
DFRQX1 DFRQX1_4 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf9), .D(_6__3_), .Q(R_3_) );
DFRQX1 DFRQX1_5 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf14), .D(_6__4_), .Q(R_4_) );
DFRQX1 DFRQX1_6 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf53), .D(_6__5_), .Q(R_5_) );
DFRQX1 DFRQX1_7 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf53), .D(_6__6_), .Q(R_6_) );
DFRQX1 DFRQX1_8 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf7), .D(_6__7_), .Q(R_7_) );
DFRQX1 DFRQX1_9 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf21), .D(_6__8_), .Q(R_8_) );
DFRQX1 DFRQX1_10 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf14), .D(_6__9_), .Q(R_9_) );
DFRQX1 DFRQX1_11 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf21), .D(_6__10_), .Q(R_10_) );
DFRQX1 DFRQX1_12 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf10), .D(_6__11_), .Q(R_11_) );
DFRQX1 DFRQX1_13 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf7), .D(_6__12_), .Q(R_12_) );
DFRQX1 DFRQX1_14 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf21), .D(_6__13_), .Q(R_13_) );
DFRQX1 DFRQX1_15 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf21), .D(_6__14_), .Q(R_14_) );
DFRQX1 DFRQX1_16 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf7), .D(_6__15_), .Q(R_15_) );
DFRQX1 DFRQX1_17 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf33), .D(_6__16_), .Q(R_16_) );
DFRQX1 DFRQX1_18 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf21), .D(_6__17_), .Q(R_17_) );
DFRQX1 DFRQX1_19 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf14), .D(_6__18_), .Q(R_18_) );
DFRQX1 DFRQX1_20 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf53), .D(_6__19_), .Q(R_19_) );
DFRQX1 DFRQX1_21 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf53), .D(_6__20_), .Q(R_20_) );
DFRQX1 DFRQX1_22 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf43), .D(_6__21_), .Q(R_21_) );
DFRQX1 DFRQX1_23 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf44), .D(_6__22_), .Q(R_22_) );
DFRQX1 DFRQX1_24 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf9), .D(_6__23_), .Q(R_23_) );
DFRQX1 DFRQX1_25 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf14), .D(_6__24_), .Q(R_24_) );
DFRQX1 DFRQX1_26 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf7), .D(_6__25_), .Q(R_25_) );
DFRQX1 DFRQX1_27 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf31), .D(_6__26_), .Q(R_26_) );
DFRQX1 DFRQX1_28 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf45), .D(_6__27_), .Q(R_27_) );
DFRQX1 DFRQX1_29 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf9), .D(_6__28_), .Q(R_28_) );
DFRQX1 DFRQX1_30 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf21), .D(_6__29_), .Q(R_29_) );
DFRQX1 DFRQX1_31 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf29), .D(_6__30_), .Q(R_30_) );
DFRQX1 DFRQX1_32 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf53), .D(_6__31_), .Q(R_31_) );
DFRQX1 DFRQX1_33 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf32), .D(_4__0_), .Q(_678__0_) );
DFRQX1 DFRQX1_34 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf23), .D(_4__1_), .Q(_678__1_) );
DFRQX1 DFRQX1_35 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf28), .D(_4__2_), .Q(_678__2_) );
DFRQX1 DFRQX1_36 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf28), .D(_4__3_), .Q(_678__3_) );
DFRQX1 DFRQX1_37 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf46), .D(_4__4_), .Q(_678__4_) );
DFRQX1 DFRQX1_38 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf23), .D(_4__5_), .Q(_678__5_) );
DFRQX1 DFRQX1_39 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf50), .D(_4__6_), .Q(_678__6_) );
DFRQX1 DFRQX1_40 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf23), .D(_4__7_), .Q(_678__7_) );
DFRQX1 DFRQX1_41 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf28), .D(_4__8_), .Q(_678__8_) );
DFRQX1 DFRQX1_42 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf23), .D(_4__9_), .Q(_678__9_) );
DFRQX1 DFRQX1_43 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf32), .D(_4__10_), .Q(_678__10_) );
DFRQX1 DFRQX1_44 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf32), .D(_4__11_), .Q(_678__11_) );
DFRQX1 DFRQX1_45 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf32), .D(_4__12_), .Q(_678__12_) );
DFRQX1 DFRQX1_46 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf28), .D(_4__13_), .Q(_678__13_) );
DFRQX1 DFRQX1_47 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf28), .D(_4__14_), .Q(_678__14_) );
DFRQX1 DFRQX1_48 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf28), .D(_4__15_), .Q(_678__15_) );
DFRQX1 DFRQX1_49 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf12), .D(_4__16_), .Q(_678__16_) );
DFRQX1 DFRQX1_50 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf32), .D(_4__17_), .Q(_678__17_) );
DFRQX1 DFRQX1_51 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf46), .D(_4__18_), .Q(_678__18_) );
DFRQX1 DFRQX1_52 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf23), .D(_4__19_), .Q(_678__19_) );
DFRQX1 DFRQX1_53 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf41), .D(_4__20_), .Q(_678__20_) );
DFRQX1 DFRQX1_54 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf23), .D(_4__21_), .Q(_678__21_) );
DFRQX1 DFRQX1_55 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf32), .D(_4__22_), .Q(_678__22_) );
DFRQX1 DFRQX1_56 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf32), .D(_4__23_), .Q(_678__23_) );
DFRQX1 DFRQX1_57 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf12), .D(_4__24_), .Q(_678__24_) );
DFRQX1 DFRQX1_58 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf50), .D(_4__25_), .Q(_678__25_) );
DFRQX1 DFRQX1_59 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf46), .D(_4__26_), .Q(_678__26_) );
DFRQX1 DFRQX1_60 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf46), .D(_4__27_), .Q(_678__27_) );
DFRQX1 DFRQX1_61 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf12), .D(_4__28_), .Q(_678__28_) );
DFRQX1 DFRQX1_62 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf28), .D(_4__29_), .Q(_678__29_) );
DFRQX1 DFRQX1_63 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf12), .D(_4__30_), .Q(_678__30_) );
DFRQX1 DFRQX1_64 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf23), .D(_4__31_), .Q(_678__31_) );
DFRQX1 DFRQX1_65 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf50), .D(_3__0_), .Q(_681__0_) );
DFRQX1 DFRQX1_66 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf1), .D(_3__1_), .Q(_681__1_) );
DFRQX1 DFRQX1_67 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf1), .D(_3__2_), .Q(_681__2_) );
DFRQX1 DFRQX1_68 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf50), .D(_3__3_), .Q(_681__3_) );
DFRQX1 DFRQX1_69 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf37), .D(_3__4_), .Q(_681__4_) );
DFRQX1 DFRQX1_70 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf1), .D(_3__5_), .Q(_681__5_) );
DFRQX1 DFRQX1_71 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf1), .D(_3__6_), .Q(_681__6_) );
DFRQX1 DFRQX1_72 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf37), .D(_3__7_), .Q(_681__7_) );
DFRQX1 DFRQX1_73 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf37), .D(_3__8_), .Q(_681__8_) );
DFRQX1 DFRQX1_74 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf27), .D(_3__9_), .Q(_681__9_) );
DFRQX1 DFRQX1_75 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf13), .D(_3__10_), .Q(_681__10_) );
DFRQX1 DFRQX1_76 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf1), .D(_3__11_), .Q(_681__11_) );
DFRQX1 DFRQX1_77 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf1), .D(_3__12_), .Q(_681__12_) );
DFRQX1 DFRQX1_78 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf37), .D(_3__13_), .Q(_681__13_) );
DFRQX1 DFRQX1_79 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf1), .D(_3__14_), .Q(_681__14_) );
DFRQX1 DFRQX1_80 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf11), .D(_3__15_), .Q(_681__15_) );
DFRQX1 DFRQX1_81 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf17), .D(_3__16_), .Q(_681__16_) );
DFRQX1 DFRQX1_82 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf37), .D(_3__17_), .Q(_681__17_) );
DFRQX1 DFRQX1_83 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf12), .D(_3__18_), .Q(_681__18_) );
DFRQX1 DFRQX1_84 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf13), .D(_3__19_), .Q(_681__19_) );
DFRQX1 DFRQX1_85 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf37), .D(_3__20_), .Q(_681__20_) );
DFRQX1 DFRQX1_86 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf37), .D(_3__21_), .Q(_681__21_) );
DFRQX1 DFRQX1_87 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf13), .D(_3__22_), .Q(_681__22_) );
DFRQX1 DFRQX1_88 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf26), .D(_3__23_), .Q(_681__23_) );
DFRQX1 DFRQX1_89 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf27), .D(_3__24_), .Q(_681__24_) );
DFRQX1 DFRQX1_90 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf12), .D(_3__25_), .Q(_681__25_) );
DFRQX1 DFRQX1_91 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf26), .D(_3__26_), .Q(_681__26_) );
DFRQX1 DFRQX1_92 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf17), .D(_3__27_), .Q(_681__27_) );
DFRQX1 DFRQX1_93 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf37), .D(_3__28_), .Q(_681__28_) );
DFRQX1 DFRQX1_94 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf11), .D(_3__29_), .Q(_681__29_) );
DFRQX1 DFRQX1_95 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf27), .D(_3__30_), .Q(_681__30_) );
DFRQX1 DFRQX1_96 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf27), .D(_3__31_), .Q(_681__31_) );
DFRQX1 DFRQX1_97 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf39), .D(_0__0_), .Q(I1_0_) );
DFRQX1 DFRQX1_98 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf42), .D(_0__1_), .Q(I1_1_) );
DFRQX1 DFRQX1_99 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf42), .D(_0__2_), .Q(I1_2_) );
DFRQX1 DFRQX1_100 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf45), .D(_0__3_), .Q(I1_3_) );
DFRQX1 DFRQX1_101 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf9), .D(_0__4_), .Q(I1_4_) );
DFRQX1 DFRQX1_102 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf29), .D(_0__5_), .Q(I1_5_) );
DFRQX1 DFRQX1_103 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf31), .D(_0__6_), .Q(I1_6_) );
DFRQX1 DFRQX1_104 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf45), .D(_0__7_), .Q(I1_7_) );
DFRQX1 DFRQX1_105 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf29), .D(_0__8_), .Q(I1_8_) );
DFRQX1 DFRQX1_106 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf8), .D(_0__9_), .Q(I1_9_) );
DFRQX1 DFRQX1_107 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf8), .D(_0__10_), .Q(I1_10_) );
DFRQX1 DFRQX1_108 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf8), .D(_0__11_), .Q(I1_11_) );
DFRQX1 DFRQX1_109 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf29), .D(_0__12_), .Q(I1_12_) );
DFRQX1 DFRQX1_110 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf4), .D(_0__13_), .Q(I1_13_) );
DFRQX1 DFRQX1_111 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf45), .D(_0__14_), .Q(I1_14_) );
DFRQX1 DFRQX1_112 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf45), .D(_0__15_), .Q(I1_15_) );
DFRQX1 DFRQX1_113 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf45), .D(_0__16_), .Q(I1_16_) );
DFRQX1 DFRQX1_114 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf42), .D(_0__17_), .Q(I1_17_) );
DFRQX1 DFRQX1_115 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf45), .D(_0__18_), .Q(I1_18_) );
DFRQX1 DFRQX1_116 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf33), .D(_0__19_), .Q(I1_19_) );
DFRQX1 DFRQX1_117 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf4), .D(_0__20_), .Q(I1_20_) );
DFRQX1 DFRQX1_118 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf4), .D(_0__21_), .Q(I1_21_) );
DFRQX1 DFRQX1_119 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf4), .D(_0__22_), .Q(I1_22_) );
DFRQX1 DFRQX1_120 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf29), .D(_0__23_), .Q(I1_23_) );
DFRQX1 DFRQX1_121 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf4), .D(_0__24_), .Q(I1_24_) );
DFRQX1 DFRQX1_122 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf8), .D(_0__25_), .Q(I1_25_) );
DFRQX1 DFRQX1_123 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf8), .D(_0__26_), .Q(I1_26_) );
DFRQX1 DFRQX1_124 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf4), .D(_0__27_), .Q(I1_27_) );
DFRQX1 DFRQX1_125 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf29), .D(_0__28_), .Q(I1_28_) );
DFRQX1 DFRQX1_126 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf45), .D(_0__29_), .Q(I1_29_) );
DFRQX1 DFRQX1_127 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf31), .D(_0__30_), .Q(I1_30_) );
DFRQX1 DFRQX1_128 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf4), .D(_0__31_), .Q(I1_31_) );
DFRRQX1 DFRRQX1_1 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf40), .D(_5__0_), .Q(_684__0_), .RN(_268__bF_buf7) );
DFRRQX1 DFRRQX1_2 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf50), .D(_5__1_), .Q(_684__1_), .RN(_268__bF_buf4) );
DFRRQX1 DFRRQX1_3 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf46), .D(_5__2_), .Q(_684__2_), .RN(_268__bF_buf7) );
DFRRQX1 DFRRQX1_4 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf50), .D(_5__3_), .Q(_684__3_), .RN(_268__bF_buf4) );
DFRRQX1 DFRRQX1_5 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf46), .D(_5__4_), .Q(_684__4_), .RN(_268__bF_buf7) );
DFRRQX1 DFRRQX1_6 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf50), .D(_5__5_), .Q(_684__5_), .RN(_268__bF_buf4) );
DFRRQX1 DFRRQX1_7 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf27), .D(_5__6_), .Q(_684__6_), .RN(_268__bF_buf8) );
DFRRQX1 DFRRQX1_8 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf31), .D(_5__7_), .Q(_684__7_), .RN(_268__bF_buf5) );
DFRRQX1 DFRRQX1_9 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf41), .D(_5__8_), .Q(_684__8_), .RN(_268__bF_buf4) );
DFRRQX1 DFRRQX1_10 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf40), .D(_5__9_), .Q(_684__9_), .RN(_268__bF_buf7) );
DFRRQX1 DFRRQX1_11 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf27), .D(_5__10_), .Q(_684__10_), .RN(_268__bF_buf8) );
DFRRQX1 DFRRQX1_12 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf40), .D(_5__11_), .Q(_684__11_), .RN(_268__bF_buf8) );
DFRRQX1 DFRRQX1_13 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf40), .D(_5__12_), .Q(_684__12_), .RN(_268__bF_buf8) );
DFRRQX1 DFRRQX1_14 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf31), .D(_5__13_), .Q(_684__13_), .RN(_268__bF_buf5) );
DFRRQX1 DFRRQX1_15 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf12), .D(_5__14_), .Q(_684__14_), .RN(_268__bF_buf7) );
DFRRQX1 DFRRQX1_16 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf26), .D(_5__15_), .Q(_684__15_), .RN(_268__bF_buf8) );
DFRRQX1 DFRRQX1_17 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf14), .D(_5__16_), .Q(_684__16_), .RN(_268__bF_buf2) );
DFRRQX1 DFRRQX1_18 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf40), .D(_5__17_), .Q(_684__17_), .RN(_268__bF_buf7) );
DFRRQX1 DFRRQX1_19 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf46), .D(_5__18_), .Q(_684__18_), .RN(_268__bF_buf7) );
DFRRQX1 DFRRQX1_20 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf40), .D(_5__19_), .Q(_684__19_), .RN(_268__bF_buf7) );
DFRRQX1 DFRRQX1_21 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf41), .D(_5__20_), .Q(_684__20_), .RN(_268__bF_buf4) );
DFRRQX1 DFRRQX1_22 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf50), .D(_5__21_), .Q(_684__21_), .RN(_268__bF_buf7) );
DFRRQX1 DFRRQX1_23 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf40), .D(_5__22_), .Q(_684__22_), .RN(_268__bF_buf8) );
DFRRQX1 DFRRQX1_24 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf40), .D(_5__23_), .Q(_684__23_), .RN(_268__bF_buf7) );
DFRRQX1 DFRRQX1_25 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf27), .D(_5__24_), .Q(_684__24_), .RN(_268__bF_buf8) );
DFRRQX1 DFRRQX1_26 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf26), .D(_5__25_), .Q(_684__25_), .RN(_268__bF_buf8) );
DFRRQX1 DFRRQX1_27 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf26), .D(_5__26_), .Q(_684__26_), .RN(_268__bF_buf8) );
DFRRQX1 DFRRQX1_28 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf14), .D(_5__27_), .Q(_684__27_), .RN(_268__bF_buf2) );
DFRRQX1 DFRRQX1_29 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf41), .D(_5__28_), .Q(_684__28_), .RN(_268__bF_buf4) );
DFRRQX1 DFRRQX1_30 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf46), .D(_5__29_), .Q(_684__29_), .RN(_268__bF_buf7) );
DFRRQX1 DFRRQX1_31 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf26), .D(_5__30_), .Q(_684__30_), .RN(_268__bF_buf8) );
DFRRQX1 DFRRQX1_32 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf26), .D(_5__31_), .Q(_684__31_), .RN(_268__bF_buf8) );
DFRRQX1 DFRRQX1_33 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf31), .D(_2__0_), .Q(PC1_0_), .RN(_268__bF_buf1) );
DFRRQX1 DFRRQX1_34 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf34), .D(_2__1_), .Q(PC1_1_), .RN(_268__bF_buf1) );
DFRRQX1 DFRRQX1_35 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf2), .D(_2__2_), .Q(PC1_2_), .RN(_268__bF_buf0) );
DFRRQX1 DFRRQX1_36 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf2), .D(_2__3_), .Q(PC1_3_), .RN(_268__bF_buf0) );
DFRRQX1 DFRRQX1_37 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf2), .D(_2__4_), .Q(PC1_4_), .RN(_268__bF_buf0) );
DFRRQX1 DFRRQX1_38 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf41), .D(_2__5_), .Q(PC1_5_), .RN(_268__bF_buf4) );
DFRRQX1 DFRRQX1_39 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf34), .D(_2__6_), .Q(PC1_6_), .RN(_268__bF_buf4) );
DFRRQX1 DFRRQX1_40 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf30), .D(_2__7_), .Q(PC1_7_), .RN(_268__bF_buf0) );
DFRRQX1 DFRRQX1_41 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf34), .D(_2__8_), .Q(PC1_8_), .RN(_268__bF_buf1) );
DFRRQX1 DFRRQX1_42 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf41), .D(_2__9_), .Q(PC1_9_), .RN(_268__bF_buf4) );
DFRRQX1 DFRRQX1_43 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf2), .D(_2__10_), .Q(PC1_10_), .RN(_268__bF_buf0) );
DFRRQX1 DFRRQX1_44 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf30), .D(_2__11_), .Q(PC1_11_), .RN(_268__bF_buf1) );
DFRRQX1 DFRRQX1_45 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf34), .D(_2__12_), .Q(PC1_12_), .RN(_268__bF_buf1) );
DFRRQX1 DFRRQX1_46 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf42), .D(_2__13_), .Q(PC1_13_), .RN(_268__bF_buf5) );
DFRRQX1 DFRRQX1_47 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf2), .D(_2__14_), .Q(PC1_14_), .RN(_268__bF_buf0) );
DFRRQX1 DFRRQX1_48 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf51), .D(_2__15_), .Q(PC1_15_), .RN(_268__bF_buf3) );
DFRRQX1 DFRRQX1_49 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf34), .D(_2__16_), .Q(PC1_16_), .RN(_268__bF_buf1) );
DFRRQX1 DFRRQX1_50 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf34), .D(_2__17_), .Q(PC1_17_), .RN(_268__bF_buf1) );
DFRRQX1 DFRRQX1_51 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf42), .D(_2__18_), .Q(PC1_18_), .RN(_268__bF_buf5) );
DFRRQX1 DFRRQX1_52 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf2), .D(_2__19_), .Q(PC1_19_), .RN(_268__bF_buf0) );
DFRRQX1 DFRRQX1_53 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf41), .D(_2__20_), .Q(PC1_20_), .RN(_268__bF_buf4) );
DFRRQX1 DFRRQX1_54 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf34), .D(_2__21_), .Q(PC1_21_), .RN(_268__bF_buf1) );
DFRRQX1 DFRRQX1_55 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf8), .D(_2__22_), .Q(PC1_22_), .RN(_268__bF_buf5) );
DFRRQX1 DFRRQX1_56 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf30), .D(_2__23_), .Q(PC1_23_), .RN(_268__bF_buf1) );
DFRRQX1 DFRRQX1_57 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf29), .D(_2__24_), .Q(PC1_24_), .RN(_268__bF_buf0) );
DFRRQX1 DFRRQX1_58 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf42), .D(_2__25_), .Q(PC1_25_), .RN(_268__bF_buf0) );
DFRRQX1 DFRRQX1_59 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf34), .D(_2__26_), .Q(PC1_26_), .RN(_268__bF_buf1) );
DFRRQX1 DFRRQX1_60 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf42), .D(_2__27_), .Q(PC1_27_), .RN(_268__bF_buf5) );
DFRRQX1 DFRRQX1_61 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf42), .D(_2__28_), .Q(PC1_28_), .RN(_268__bF_buf5) );
DFRRQX1 DFRRQX1_62 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf2), .D(_2__29_), .Q(PC1_29_), .RN(_268__bF_buf0) );
DFRRQX1 DFRRQX1_63 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf31), .D(_2__30_), .Q(PC1_30_), .RN(_268__bF_buf5) );
DFRRQX1 DFRRQX1_64 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf9), .D(_2__31_), .Q(PC1_31_), .RN(_268__bF_buf5) );
DFRSQX1 DFRSQX1_1 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf53), .D(_1__0_), .Q(CTRL_IDEC0_IR_0_), .SN(_268__bF_buf2) );
DFRSQX1 DFRSQX1_2 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf53), .D(_1__1_), .Q(CTRL_IDEC0_IR_1_), .SN(_268__bF_buf2) );
DFRRQX2 DFRRQX2_1 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf43), .D(_1__2_), .Q(CTRL_IDEC0_IR_2_), .RN(_268__bF_buf3) );
DFRRQX2 DFRRQX2_2 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf43), .D(_1__3_), .Q(CTRL_IDEC0_IR_3_), .RN(_268__bF_buf2) );
DFRSQX1 DFRSQX1_3 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf43), .D(_1__4_), .Q(CTRL_IDEC0_IR_4_), .SN(_268__bF_buf3) );
DFRRQX1 DFRRQX1_65 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf41), .D(_1__5_), .Q(CTRL_IDEC0_IR_5_), .RN(_268__bF_buf4) );
DFRRQX2 DFRRQX2_3 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf9), .D(_1__6_), .Q(CTRL_IDEC0_IR_6_), .RN(_268__bF_buf3) );
DFRRQX1 DFRRQX1_66 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf44), .D(_1__7_), .Q(CTRL_IDEC0_IR_7_), .RN(_268__bF_buf6) );
DFRRQX1 DFRRQX1_67 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf8), .D(_1__8_), .Q(CTRL_IDEC0_IR_8_), .RN(_268__bF_buf5) );
DFRRQX1 DFRRQX1_68 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf44), .D(_1__9_), .Q(CTRL_IDEC0_IR_9_), .RN(_268__bF_buf2) );
DFRRQX1 DFRRQX1_69 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf33), .D(_1__10_), .Q(CTRL_IDEC0_IR_10_), .RN(_268__bF_buf3) );
DFRRQX1 DFRRQX1_70 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf0), .D(_1__11_), .Q(CTRL_IDEC0_IR_11_), .RN(_268__bF_buf3) );
DFRRQX1 DFRRQX1_71 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf39), .D(_1__12_), .Q(CTRL_IDEC0_IR_12_), .RN(_268__bF_buf6) );
DFRRQX1 DFRRQX1_72 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf44), .D(_1__13_), .Q(CTRL_IDEC0_IR_13_), .RN(_268__bF_buf6) );
DFRRQX1 DFRRQX1_73 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf43), .D(_1__14_), .Q(CTRL_IDEC0_IR_14_), .RN(_268__bF_buf2) );
DFRRQX1 DFRRQX1_74 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf39), .D(_1__15_), .Q(_686__0_), .RN(_268__bF_buf6) );
DFRRQX1 DFRRQX1_75 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf24), .D(_1__16_), .Q(_686__1_), .RN(_268__bF_buf6) );
DFRRQX1 DFRRQX1_76 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf7), .D(_1__17_), .Q(_686__2_), .RN(_268__bF_buf2) );
DFRRQX1 DFRRQX1_77 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf43), .D(_1__18_), .Q(_686__3_), .RN(_268__bF_buf2) );
DFRRQX1 DFRRQX1_78 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf44), .D(_1__19_), .Q(_686__4_), .RN(_268__bF_buf2) );
DFRRQX2 DFRRQX2_4 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf24), .D(_1__20_), .Q(_687__0_), .RN(_268__bF_buf6) );
DFRRQX1 DFRRQX1_79 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf39), .D(_1__21_), .Q(_687__1_), .RN(_268__bF_buf6) );
DFRRQX1 DFRRQX1_80 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf24), .D(_1__22_), .Q(_687__2_), .RN(_268__bF_buf6) );
DFRRQX1 DFRRQX1_81 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf24), .D(_1__23_), .Q(_687__3_), .RN(_268__bF_buf6) );
DFRRQX1 DFRRQX1_82 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf44), .D(_1__24_), .Q(_687__4_), .RN(_268__bF_buf6) );
DFRRQX1 DFRRQX1_83 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf39), .D(_1__25_), .Q(CTRL_IDEC0_IR_25_), .RN(_268__bF_buf3) );
DFRRQX1 DFRRQX1_84 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf9), .D(_1__26_), .Q(CTRL_IDEC0_IR_26_), .RN(_268__bF_buf5) );
DFRRQX1 DFRRQX1_85 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf39), .D(_1__27_), .Q(CTRL_IDEC0_IR_27_), .RN(_268__bF_buf3) );
DFRRQX1 DFRRQX1_86 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf43), .D(_1__28_), .Q(CTRL_IDEC0_IR_28_), .RN(_268__bF_buf3) );
DFRRQX1 DFRRQX1_87 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf39), .D(_1__29_), .Q(CTRL_IDEC0_IR_29_), .RN(_268__bF_buf3) );
DFRRQX1 DFRRQX1_88 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf43), .D(_1__30_), .Q(CTRL_IDEC0_IR_30_), .RN(_268__bF_buf3) );
DFRRQX1 DFRRQX1_89 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf24), .D(_1__31_), .Q(CTRL_IDEC0_IR_31_), .RN(_268__bF_buf6) );
INX1 INX1_67 ( .gnd!(gnd!), .vdd!(vdd!), .A(_682__0_bF_buf0), .Q(_834_) );
NO2X1 NO2X1_96 ( .gnd!(gnd!), .vdd!(vdd!), .A(_682__1_bF_buf1), .B(_834_), .Q(_855_) );
INX1 INX1_68 ( .gnd!(gnd!), .vdd!(vdd!), .A(_855_), .Q(_856_) );
INX2 INX2_5 ( .gnd!(gnd!), .vdd!(vdd!), .A(EXT_type_bF_buf2), .Q(_866_) );
NO2X1 NO2X1_97 ( .gnd!(gnd!), .vdd!(vdd!), .A(ALU_opcode_1_), .B(ALU_opcode_0_), .Q(_877_) );
NA3I1X2 NA3I1X2_3 ( .gnd!(gnd!), .vdd!(vdd!), .AN(ALU_opcode_4_), .B(ALU_opcode_2_), .C(_877_), .Q(_888_) );
NO2X1 NO2X1_98 ( .gnd!(gnd!), .vdd!(vdd!), .A(_866__bF_buf3), .B(_888__bF_buf4), .Q(_898_) );
NA2X2 NA2X2_1 ( .gnd!(gnd!), .vdd!(vdd!), .A(_856_), .B(_898_), .Q(_909_) );
INX1 INX1_69 ( .gnd!(gnd!), .vdd!(vdd!), .A(_682__1_bF_buf1), .Q(_920_) );
NO3X2 NO3X2_1 ( .gnd!(gnd!), .vdd!(vdd!), .A(_888__bF_buf4), .B(EXT_type_bF_buf3), .C(_920_), .Q(_931_) );
NO2X2 NO2X2_1 ( .gnd!(gnd!), .vdd!(vdd!), .A(_888__bF_buf4), .B(_856_), .Q(_941_) );
INX2 INX2_6 ( .gnd!(gnd!), .vdd!(vdd!), .A(_941__bF_buf0), .Q(_952_) );
INX1 INX1_70 ( .gnd!(gnd!), .vdd!(vdd!), .A(ALU_a_0_), .Q(_963_) );
INX1 INX1_71 ( .gnd!(gnd!), .vdd!(vdd!), .A(ALU_b_0_), .Q(_973_) );
NO2X1 NO2X1_99 ( .gnd!(gnd!), .vdd!(vdd!), .A(_963_), .B(_973_), .Q(_984_) );
INX1 INX1_72 ( .gnd!(gnd!), .vdd!(vdd!), .A(_984_), .Q(_995_) );
INX1 INX1_73 ( .gnd!(gnd!), .vdd!(vdd!), .A(ALU_opcode_3_), .Q(_1005_) );
NA2I1X1 NA2I1X1_34 ( .gnd!(gnd!), .vdd!(vdd!), .AN(EXT_type_bF_buf0), .B(ALU_func7_5_bF_buf3), .Q(_1016_) );
NA3I2X1 NA3I2X1_1 ( .gnd!(gnd!), .vdd!(vdd!), .AN(_682__0_bF_buf2), .BN(_682__1_bF_buf4), .C(ALU_opcode_3_), .Q(_1027_) );
NA3I1X1 NA3I1X1_1 ( .gnd!(gnd!), .vdd!(vdd!), .AN(ALU_opcode_2_), .B(ALU_opcode_4_), .C(_877_), .Q(_1037_) );
ON32X2 ON32X2_1 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1016_), .B(_1027_), .C(_888__bF_buf0), .D(_1005_), .E(_1037_), .Q(_1048_) );
NO2X1 NO2X1_100 ( .gnd!(gnd!), .vdd!(vdd!), .A(_931__bF_buf2), .B(_1048__bF_buf4), .Q(_1059_) );
ON21X1 ON21X1_181 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1059__bF_buf2), .B(ALU_b_0_), .C(_995_), .Q(_1069_) );
INX1 INX1_74 ( .gnd!(gnd!), .vdd!(vdd!), .A(ALU_a_1_), .Q(_1080_) );
ON21X1 ON21X1_182 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1048__bF_buf4), .B(_931__bF_buf2), .C(ALU_b_1_), .Q(_1091_) );
NO2I1X1 NO2I1X1_33 ( .gnd!(gnd!), .vdd!(vdd!), .AN(ALU_opcode_2_), .B(ALU_opcode_4_), .Q(_1101_) );
NO3I1X1 NO3I1X1_1 ( .gnd!(gnd!), .vdd!(vdd!), .AN(_682__1_bF_buf1), .B(EXT_type_bF_buf3), .C(_682__0_bF_buf0), .Q(_1112_) );
NA2X1 NA2X1_168 ( .gnd!(gnd!), .vdd!(vdd!), .A(_682__0_bF_buf2), .B(_682__1_bF_buf4), .Q(_1123_) );
NO2X1 NO2X1_101 ( .gnd!(gnd!), .vdd!(vdd!), .A(EXT_type_bF_buf3), .B(_1123_), .Q(_1133_) );
ON211X2 ON211X2_1 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1112_), .B(_1133_), .C(_1101_), .D(_877_), .Q(_1143_) );
NA2I1X1 NA2I1X1_35 ( .gnd!(gnd!), .vdd!(vdd!), .AN(ALU_opcode_4_), .B(ALU_opcode_2_), .Q(_1154_) );
NO3X1 NO3X1_1 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1154_), .B(ALU_opcode_1_), .C(ALU_opcode_0_), .Q(_1163_) );
NO2X1 NO2X1_102 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1016_), .B(_1027_), .Q(_1174_) );
NA2X1 NA2X1_169 ( .gnd!(gnd!), .vdd!(vdd!), .A(ALU_opcode_4_), .B(ALU_opcode_3_), .Q(_1185_) );
NO2X1 NO2X1_103 ( .gnd!(gnd!), .vdd!(vdd!), .A(ALU_opcode_2_), .B(_1185_), .Q(_1194_) );
AN22X2 AN22X2_1 ( .gnd!(gnd!), .vdd!(vdd!), .A(_877_), .B(_1194_), .C(_1174_), .D(_1163_), .Q(_1203_) );
NA3I1X1 NA3I1X1_2 ( .gnd!(gnd!), .vdd!(vdd!), .AN(ALU_b_1_), .B(_1143__bF_buf1), .C(_1203__bF_buf0), .Q(_1204_) );
NA3I1X1 NA3I1X1_3 ( .gnd!(gnd!), .vdd!(vdd!), .AN(_1080_), .B(_1091_), .C(_1204_), .Q(_1205_) );
INX1 INX1_75 ( .gnd!(gnd!), .vdd!(vdd!), .A(ALU_b_1_), .Q(_1206_) );
ON21X1 ON21X1_183 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1048__bF_buf4), .B(_931__bF_buf3), .C(_1206_), .Q(_1207_) );
NA3I1X1 NA3I1X1_4 ( .gnd!(gnd!), .vdd!(vdd!), .AN(_1206_), .B(_1143__bF_buf1), .C(_1203__bF_buf0), .Q(_1208_) );
NA3I1X1 NA3I1X1_5 ( .gnd!(gnd!), .vdd!(vdd!), .AN(ALU_a_1_), .B(_1207_), .C(_1208_), .Q(_1209_) );
NA3X1 NA3X1_1 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1069_), .B(_1205_), .C(_1209_), .Q(_1210_) );
NA2X1 NA2X1_170 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1194_), .B(_877_), .Q(_1211_) );
ON311X2 ON311X2_1 ( .gnd!(gnd!), .vdd!(vdd!), .A(_888__bF_buf3), .B(_1016_), .C(_1027_), .D(_1211_), .E(_1143__bF_buf1), .Q(_1212_) );
AN21X1 AN21X1_77 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1212__bF_buf3), .B(_973_), .C(_984_), .Q(_1213_) );
NA3I1X1 NA3I1X1_6 ( .gnd!(gnd!), .vdd!(vdd!), .AN(ALU_a_1_), .B(_1091_), .C(_1204_), .Q(_1214_) );
NA3I1X1 NA3I1X1_7 ( .gnd!(gnd!), .vdd!(vdd!), .AN(_1080_), .B(_1207_), .C(_1208_), .Q(_1215_) );
NA3X1 NA3X1_2 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1213_), .B(_1214_), .C(_1215_), .Q(_1216_) );
NA2X1 NA2X1_171 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1163_), .B(_1005_), .Q(_1217_) );
NA2X1 NA2X1_172 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1217_), .B(ALU_b_4_), .Q(_1218_) );
NO2X1 NO2X1_104 ( .gnd!(gnd!), .vdd!(vdd!), .A(ALU_opcode_3_), .B(_888__bF_buf4), .Q(_1219_) );
NA2X1 NA2X1_173 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1219_), .B(ALU_shamt_4_), .Q(_1220_) );
NA2X2 NA2X2_2 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1218_), .B(_1220_), .Q(_1221_) );
INX2 INX2_7 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1221__bF_buf1), .Q(_1222_) );
INX1 INX1_76 ( .gnd!(gnd!), .vdd!(vdd!), .A(ALU_func7_5_bF_buf2), .Q(_1223_) );
NA2X1 NA2X1_174 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1217_), .B(ALU_b_3_), .Q(_1224_) );
NA2X1 NA2X1_175 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1219_), .B(ALU_shamt_3_), .Q(_1225_) );
NA2X3 NA2X3_1 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1224_), .B(_1225_), .Q(_1226_) );
INX3 INX3_6 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1226__bF_buf1), .Q(_1227_) );
NA2X1 NA2X1_176 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1217_), .B(ALU_b_2_), .Q(_1228_) );
NA2X1 NA2X1_177 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1219_), .B(ALU_shamt_2_), .Q(_1229_) );
NA2X3 NA2X3_2 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1228_), .B(_1229_), .Q(_1230_) );
NA2X1 NA2X1_178 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1217_), .B(ALU_b_1_), .Q(_1231_) );
NA2X1 NA2X1_179 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1219_), .B(ALU_shamt_1_), .Q(_1232_) );
AND2X2 AND2X2_2 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1231_), .B(_1232_), .Q(_1233_) );
NA2X1 NA2X1_180 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1219_), .B(CTRL_cu_csr_rd_s1_bF_buf5), .Q(_1234_) );
ON21X2 ON21X2_1 ( .gnd!(gnd!), .vdd!(vdd!), .A(_973_), .B(_1219_), .C(_1234_), .Q(_1235_) );
MU2IX1 MU2IX1_13 ( .gnd!(gnd!), .vdd!(vdd!), .IN0(ALU_a_23_), .IN1(ALU_a_24_), .Q(_1236_), .S(_1235__bF_buf4) );
MU2IX1 MU2IX1_14 ( .gnd!(gnd!), .vdd!(vdd!), .IN0(ALU_a_21_), .IN1(ALU_a_22_), .Q(_1237_), .S(_1235__bF_buf4) );
MU2IX1 MU2IX1_15 ( .gnd!(gnd!), .vdd!(vdd!), .IN0(_1236_), .IN1(_1237_), .Q(_1238_), .S(_1233__bF_buf2) );
NA2X1 NA2X1_181 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1238_), .B(_1230__bF_buf4), .Q(_1239_) );
NA2X3 NA2X3_3 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1231_), .B(_1232_), .Q(_1240_) );
NA2I1X1 NA2I1X1_36 ( .gnd!(gnd!), .vdd!(vdd!), .AN(CTRL_cu_csr_rd_s1_bF_buf5), .B(_1219_), .Q(_1241_) );
ON21X2 ON21X2_2 ( .gnd!(gnd!), .vdd!(vdd!), .A(ALU_b_0_), .B(_1219_), .C(_1241_), .Q(_1242_) );
NA2X1 NA2X1_182 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1242__bF_buf0), .B(ALU_a_19_), .Q(_1243_) );
NA2X1 NA2X1_183 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1235__bF_buf3), .B(ALU_a_20_), .Q(_1244_) );
AND2X2 AND2X2_3 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1243_), .B(_1244_), .Q(_1245_) );
NA2X1 NA2X1_184 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1242__bF_buf0), .B(ALU_a_17_), .Q(_1246_) );
NA2X1 NA2X1_185 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1235__bF_buf3), .B(ALU_a_18_), .Q(_1247_) );
NA2X1 NA2X1_186 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1246_), .B(_1247_), .Q(_1248_) );
INX1 INX1_77 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1248_), .Q(_1249_) );
MU2X1 MU2X1_170 ( .gnd!(gnd!), .vdd!(vdd!), .IN0(_1249_), .IN1(_1245_), .Q(_1250_), .S(_1240__bF_buf1) );
ON211X1 ON211X1_34 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1250_), .B(_1230__bF_buf4), .C(_1227__bF_buf4), .D(_1239_), .Q(_1251_) );
INX3 INX3_7 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1230__bF_buf0), .Q(_1252_) );
MU2IX1 MU2IX1_16 ( .gnd!(gnd!), .vdd!(vdd!), .IN0(ALU_a_27_), .IN1(ALU_a_28_), .Q(_1253_), .S(_1235__bF_buf1) );
MU2IX1 MU2IX1_17 ( .gnd!(gnd!), .vdd!(vdd!), .IN0(ALU_a_25_), .IN1(ALU_a_26_), .Q(_1254_), .S(_1235__bF_buf1) );
MU2IX1 MU2IX1_18 ( .gnd!(gnd!), .vdd!(vdd!), .IN0(_1253_), .IN1(_1254_), .Q(_1255_), .S(_1233__bF_buf2) );
NA2X1 NA2X1_187 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1242__bF_buf1), .B(ALU_a_29_), .Q(_1256_) );
NA2X1 NA2X1_188 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1235__bF_buf4), .B(ALU_a_30_), .Q(_1257_) );
AND2X2 AND2X2_4 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1256_), .B(_1257_), .Q(_1258_) );
NA2X1 NA2X1_189 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1240__bF_buf1), .B(ALU_a_31_), .Q(_1259_) );
ON21X1 ON21X1_184 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1258_), .B(_1240__bF_buf1), .C(_1259_), .Q(_1260_) );
MU2X1 MU2X1_171 ( .gnd!(gnd!), .vdd!(vdd!), .IN0(_1260_), .IN1(_1255_), .Q(_1261_), .S(_1252__bF_buf5) );
ON21X1 ON21X1_185 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1227__bF_buf2), .B(_1261_), .C(_1251_), .Q(_1262_) );
NA2I1X1 NA2I1X1_37 ( .gnd!(gnd!), .vdd!(vdd!), .AN(_1255_), .B(_1252__bF_buf5), .Q(_1263_) );
NA2X1 NA2X1_190 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1256_), .B(_1257_), .Q(_1264_) );
INX1 INX1_78 ( .gnd!(gnd!), .vdd!(vdd!), .A(ALU_a_31_), .Q(_1265_) );
NO2X1 NO2X1_105 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1265_), .B(_1235__bF_buf1), .Q(_1266_) );
MU2IX1 MU2IX1_19 ( .gnd!(gnd!), .vdd!(vdd!), .IN0(_1264_), .IN1(_1266_), .Q(_1267_), .S(_1240__bF_buf1) );
NA2X1 NA2X1_191 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1267_), .B(_1230__bF_buf4), .Q(_1268_) );
NA2X1 NA2X1_192 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1263_), .B(_1268_), .Q(_1269_) );
NA2X1 NA2X1_193 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1269_), .B(_1226__bF_buf4), .Q(_1270_) );
NA2X1 NA2X1_194 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1270_), .B(_1251_), .Q(_1271_) );
MU2IX1 MU2IX1_20 ( .gnd!(gnd!), .vdd!(vdd!), .IN0(_1262_), .IN1(_1271_), .Q(_1272_), .S(_1223_) );
INX1 INX1_79 ( .gnd!(gnd!), .vdd!(vdd!), .A(ALU_a_15_), .Q(_1273_) );
NA2X1 NA2X1_195 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1242__bF_buf2), .B(_1273_), .Q(_1274_) );
ON21X1 ON21X1_186 ( .gnd!(gnd!), .vdd!(vdd!), .A(ALU_a_16_), .B(_1242__bF_buf0), .C(_1274_), .Q(_1275_) );
INX1 INX1_80 ( .gnd!(gnd!), .vdd!(vdd!), .A(ALU_a_13_), .Q(_1276_) );
NA2X1 NA2X1_196 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1242__bF_buf2), .B(_1276_), .Q(_1277_) );
INX1 INX1_81 ( .gnd!(gnd!), .vdd!(vdd!), .A(ALU_a_14_), .Q(_1278_) );
NA2X1 NA2X1_197 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1235__bF_buf2), .B(_1278_), .Q(_1279_) );
NA2X1 NA2X1_198 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1277_), .B(_1279_), .Q(_1280_) );
MU2IX1 MU2IX1_21 ( .gnd!(gnd!), .vdd!(vdd!), .IN0(_1280_), .IN1(_1275_), .Q(_1281_), .S(_1240__bF_buf5) );
INX1 INX1_82 ( .gnd!(gnd!), .vdd!(vdd!), .A(ALU_a_11_), .Q(_1282_) );
NA2X1 NA2X1_199 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1242__bF_buf2), .B(_1282_), .Q(_1283_) );
INX1 INX1_83 ( .gnd!(gnd!), .vdd!(vdd!), .A(ALU_a_12_), .Q(_1284_) );
NA2X1 NA2X1_200 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1235__bF_buf2), .B(_1284_), .Q(_1285_) );
NA2X1 NA2X1_201 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1283_), .B(_1285_), .Q(_1286_) );
INX1 INX1_84 ( .gnd!(gnd!), .vdd!(vdd!), .A(ALU_a_9_), .Q(_1287_) );
NA2X1 NA2X1_202 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1242__bF_buf4), .B(_1287_), .Q(_1288_) );
INX1 INX1_85 ( .gnd!(gnd!), .vdd!(vdd!), .A(ALU_a_10_), .Q(_1289_) );
NA2X1 NA2X1_203 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1235__bF_buf2), .B(_1289_), .Q(_1290_) );
NA2X1 NA2X1_204 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1288_), .B(_1290_), .Q(_1291_) );
MU2IX1 MU2IX1_22 ( .gnd!(gnd!), .vdd!(vdd!), .IN0(_1291_), .IN1(_1286_), .Q(_1292_), .S(_1240__bF_buf5) );
MU2X1 MU2X1_172 ( .gnd!(gnd!), .vdd!(vdd!), .IN0(_1281_), .IN1(_1292_), .Q(_1293_), .S(_1252__bF_buf5) );
NA2X1 NA2X1_205 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1293_), .B(_1226__bF_buf1), .Q(_1294_) );
INX1 INX1_86 ( .gnd!(gnd!), .vdd!(vdd!), .A(ALU_a_3_), .Q(_1295_) );
NA2X1 NA2X1_206 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1242__bF_buf4), .B(_1295_), .Q(_1296_) );
INX1 INX1_87 ( .gnd!(gnd!), .vdd!(vdd!), .A(ALU_a_4_), .Q(_1297_) );
NA2X1 NA2X1_207 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1235__bF_buf0), .B(_1297_), .Q(_1298_) );
NA2X1 NA2X1_208 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1296_), .B(_1298_), .Q(_1299_) );
NO2X1 NO2X1_106 ( .gnd!(gnd!), .vdd!(vdd!), .A(ALU_a_2_), .B(_1242__bF_buf3), .Q(_1300_) );
NA2X1 NA2X1_209 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1242__bF_buf3), .B(_1080_), .Q(_1301_) );
NA2X1 NA2X1_210 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1233__bF_buf0), .B(_1301_), .Q(_1302_) );
ON22X1 ON22X1_1 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1302_), .B(_1300_), .C(_1299_), .D(_1233__bF_buf0), .Q(_1303_) );
INX1 INX1_88 ( .gnd!(gnd!), .vdd!(vdd!), .A(ALU_a_7_), .Q(_1304_) );
NA2X1 NA2X1_211 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1242__bF_buf4), .B(_1304_), .Q(_1305_) );
INX1 INX1_89 ( .gnd!(gnd!), .vdd!(vdd!), .A(ALU_a_8_), .Q(_1306_) );
NA2X1 NA2X1_212 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1235__bF_buf2), .B(_1306_), .Q(_1307_) );
NA2X1 NA2X1_213 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1305_), .B(_1307_), .Q(_1308_) );
INX1 INX1_90 ( .gnd!(gnd!), .vdd!(vdd!), .A(ALU_a_5_), .Q(_1309_) );
NA2X1 NA2X1_214 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1242__bF_buf4), .B(_1309_), .Q(_1310_) );
INX1 INX1_91 ( .gnd!(gnd!), .vdd!(vdd!), .A(ALU_a_6_), .Q(_1311_) );
NA2X1 NA2X1_215 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1235__bF_buf0), .B(_1311_), .Q(_1312_) );
NA2X1 NA2X1_216 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1310_), .B(_1312_), .Q(_1313_) );
MU2IX1 MU2IX1_23 ( .gnd!(gnd!), .vdd!(vdd!), .IN0(_1313_), .IN1(_1308_), .Q(_1314_), .S(_1240__bF_buf3) );
MU2IX1 MU2IX1_24 ( .gnd!(gnd!), .vdd!(vdd!), .IN0(_1303_), .IN1(_1314_), .Q(_1315_), .S(_1230__bF_buf3) );
ON211X1 ON211X1_35 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1226__bF_buf1), .B(_1315_), .C(_1294_), .D(_1222__bF_buf5), .Q(_1316_) );
ON211X1 ON211X1_36 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1272_), .B(_1222__bF_buf5), .C(EXT_type_bF_buf4), .D(_1316_), .Q(_1317_) );
ON21X1 ON21X1_187 ( .gnd!(gnd!), .vdd!(vdd!), .A(ALU_a_0_), .B(_1242__bF_buf3), .C(_1301_), .Q(_1318_) );
NO2X1 NO2X1_107 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1240__bF_buf0), .B(_1318_), .Q(_1319_) );
NA2X1 NA2X1_217 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1319_), .B(_1252__bF_buf4), .Q(_1320_) );
NO2X1 NO2X1_108 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1226__bF_buf5), .B(_1320_), .Q(_1321_) );
NO2X1 NO2X1_109 ( .gnd!(gnd!), .vdd!(vdd!), .A(EXT_type_bF_buf6), .B(_1221__bF_buf0), .Q(_1322_) );
NA2X1 NA2X1_218 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1321_), .B(_1322__bF_buf1), .Q(_1323_) );
AN21X1 AN21X1_78 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1317_), .B(_1323_), .C(_952__bF_buf0), .Q(_1324_) );
AN31X1 AN31X1_33 ( .gnd!(gnd!), .vdd!(vdd!), .A(_952__bF_buf4), .B(_1210_), .C(_1216_), .D(_1324_), .Q(_1325_) );
NO3X1 NO3X1_2 ( .gnd!(gnd!), .vdd!(vdd!), .A(_866__bF_buf5), .B(_920_), .C(_682__0_bF_buf0), .Q(_1326_) );
NA2X1 NA2X1_219 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1326_), .B(_1163_), .Q(_1327_) );
INX2 INX2_8 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1327_), .Q(_1328_) );
NA2I1X2 NA2I1X2_1 ( .gnd!(gnd!), .vdd!(vdd!), .AN(_1123_), .B(EXT_type_bF_buf3), .Q(_1329_) );
NO2X1 NO2X1_110 ( .gnd!(gnd!), .vdd!(vdd!), .A(_888__bF_buf3), .B(_1329__bF_buf0), .Q(_1330_) );
AN21X1 AN21X1_79 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1080_), .B(_1206_), .C(_1330_), .Q(_1331_) );
ON31X1 ON31X1_33 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1080_), .B(_1206_), .C(_1328__bF_buf0), .D(_1331_), .Q(_1332_) );
AN31X1 AN31X1_34 ( .gnd!(gnd!), .vdd!(vdd!), .A(ALU_a_1_), .B(ALU_b_1_), .C(_1330_), .D(_909__bF_buf2), .Q(_1333_) );
AN221X1 AN221X1_1 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1332_), .B(_1333_), .C(_1325_), .D(_909__bF_buf0), .E(_931__bF_buf3), .Q(ALU_r_1_) );
NA2X1 NA2X1_220 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1242__bF_buf1), .B(ALU_a_24_), .Q(_1334_) );
NA2X1 NA2X1_221 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1235__bF_buf1), .B(ALU_a_25_), .Q(_1335_) );
NA2X1 NA2X1_222 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1334_), .B(_1335_), .Q(_1336_) );
NA2X1 NA2X1_223 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1242__bF_buf1), .B(ALU_a_22_), .Q(_1337_) );
NA2X1 NA2X1_224 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1235__bF_buf4), .B(ALU_a_23_), .Q(_1338_) );
NA2X1 NA2X1_225 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1337_), .B(_1338_), .Q(_1339_) );
MU2X1 MU2X1_173 ( .gnd!(gnd!), .vdd!(vdd!), .IN0(_1339_), .IN1(_1336_), .Q(_1340_), .S(_1240__bF_buf5) );
NA2X1 NA2X1_226 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1242__bF_buf0), .B(ALU_a_20_), .Q(_1341_) );
NA2X1 NA2X1_227 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1235__bF_buf3), .B(ALU_a_21_), .Q(_1342_) );
NA2X1 NA2X1_228 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1341_), .B(_1342_), .Q(_1343_) );
NA2X1 NA2X1_229 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1242__bF_buf0), .B(ALU_a_18_), .Q(_1344_) );
NA2X1 NA2X1_230 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1235__bF_buf3), .B(ALU_a_19_), .Q(_1345_) );
NA2X1 NA2X1_231 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1344_), .B(_1345_), .Q(_1346_) );
MU2X1 MU2X1_174 ( .gnd!(gnd!), .vdd!(vdd!), .IN0(_1346_), .IN1(_1343_), .Q(_1347_), .S(_1240__bF_buf4) );
MU2X1 MU2X1_175 ( .gnd!(gnd!), .vdd!(vdd!), .IN0(_1347_), .IN1(_1340_), .Q(_1348_), .S(_1230__bF_buf5) );
NA2X1 NA2X1_232 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1242__bF_buf1), .B(ALU_a_28_), .Q(_1349_) );
NA2X1 NA2X1_233 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1235__bF_buf1), .B(ALU_a_29_), .Q(_1350_) );
NA2X1 NA2X1_234 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1349_), .B(_1350_), .Q(_1351_) );
NA2X1 NA2X1_235 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1351_), .B(_1240__bF_buf1), .Q(_1352_) );
NA2X1 NA2X1_236 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1242__bF_buf1), .B(ALU_a_26_), .Q(_1353_) );
NA2X1 NA2X1_237 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1235__bF_buf1), .B(ALU_a_27_), .Q(_1354_) );
NA2X1 NA2X1_238 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1353_), .B(_1354_), .Q(_1355_) );
NA2X1 NA2X1_239 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1355_), .B(_1233__bF_buf1), .Q(_1356_) );
NA2X1 NA2X1_240 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1352_), .B(_1356_), .Q(_1357_) );
NO2X1 NO2X1_111 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1230__bF_buf5), .B(_1357_), .Q(_1358_) );
NA2X1 NA2X1_241 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1242__bF_buf1), .B(ALU_a_30_), .Q(_1359_) );
ON21X1 ON21X1_188 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1265_), .B(_1242__bF_buf1), .C(_1359_), .Q(_1360_) );
NA2X1 NA2X1_242 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1360_), .B(_1233__bF_buf1), .Q(_1361_) );
AN21X1 AN21X1_80 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1230__bF_buf5), .B(_1361_), .C(_1358_), .Q(_1362_) );
MU2X1 MU2X1_176 ( .gnd!(gnd!), .vdd!(vdd!), .IN0(_1348_), .IN1(_1362_), .Q(_1363_), .S(_1226__bF_buf3) );
NA2X1 NA2X1_243 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1363_), .B(_1223_), .Q(_1364_) );
AN31X1 AN31X1_35 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1230__bF_buf5), .B(_1259_), .C(_1361_), .D(_1358_), .Q(_1365_) );
MU2IX1 MU2IX1_25 ( .gnd!(gnd!), .vdd!(vdd!), .IN0(_1365_), .IN1(_1348_), .Q(_1366_), .S(_1227__bF_buf1) );
NA2I1X1 NA2I1X1_38 ( .gnd!(gnd!), .vdd!(vdd!), .AN(_1366_), .B(ALU_func7_5_bF_buf1), .Q(_1367_) );
NA2X1 NA2X1_244 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1242__bF_buf4), .B(_1297_), .Q(_1368_) );
NA2X1 NA2X1_245 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1235__bF_buf0), .B(_1309_), .Q(_1369_) );
AND2X2 AND2X2_5 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1368_), .B(_1369_), .Q(_1370_) );
NA2X1 NA2X1_246 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1242__bF_buf3), .B(ALU_a_2_), .Q(_1371_) );
ON21X1 ON21X1_189 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1295_), .B(_1242__bF_buf3), .C(_1371_), .Q(_1372_) );
MU2IX1 MU2IX1_26 ( .gnd!(gnd!), .vdd!(vdd!), .IN0(_1370_), .IN1(_1372_), .Q(_1373_), .S(_1233__bF_buf0) );
NA2X1 NA2X1_247 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1242__bF_buf4), .B(_1306_), .Q(_1374_) );
NA2X1 NA2X1_248 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1235__bF_buf2), .B(_1287_), .Q(_1375_) );
NA2X1 NA2X1_249 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1374_), .B(_1375_), .Q(_1376_) );
NA2X1 NA2X1_250 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1242__bF_buf4), .B(_1311_), .Q(_1377_) );
NA2X1 NA2X1_251 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1235__bF_buf0), .B(_1304_), .Q(_1378_) );
NA2X1 NA2X1_252 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1377_), .B(_1378_), .Q(_1379_) );
MU2IX1 MU2IX1_27 ( .gnd!(gnd!), .vdd!(vdd!), .IN0(_1379_), .IN1(_1376_), .Q(_1380_), .S(_1240__bF_buf6) );
NO2X1 NO2X1_112 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1252__bF_buf3), .B(_1380_), .Q(_1381_) );
AN211X1 AN211X1_1 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1252__bF_buf3), .B(_1373_), .C(_1226__bF_buf2), .D(_1381_), .Q(_1382_) );
NA2X1 NA2X1_253 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1242__bF_buf0), .B(ALU_a_16_), .Q(_1383_) );
NA2X1 NA2X1_254 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1235__bF_buf3), .B(ALU_a_17_), .Q(_1384_) );
NA2X1 NA2X1_255 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1383_), .B(_1384_), .Q(_1385_) );
NA2X1 NA2X1_256 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1385_), .B(_1240__bF_buf4), .Q(_1386_) );
NA2X1 NA2X1_257 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1242__bF_buf2), .B(_1278_), .Q(_1387_) );
ON21X1 ON21X1_190 ( .gnd!(gnd!), .vdd!(vdd!), .A(ALU_a_15_), .B(_1242__bF_buf2), .C(_1387_), .Q(_1388_) );
ON21X1 ON21X1_191 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1240__bF_buf4), .B(_1388_), .C(_1386_), .Q(_1389_) );
NA2X1 NA2X1_258 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1242__bF_buf2), .B(_1284_), .Q(_1390_) );
NA2X1 NA2X1_259 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1235__bF_buf3), .B(_1276_), .Q(_1391_) );
NA2X1 NA2X1_260 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1390_), .B(_1391_), .Q(_1392_) );
NA2X1 NA2X1_261 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1242__bF_buf2), .B(_1289_), .Q(_1393_) );
NA2X1 NA2X1_262 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1235__bF_buf2), .B(_1282_), .Q(_1394_) );
NA2X1 NA2X1_263 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1393_), .B(_1394_), .Q(_1395_) );
MU2IX1 MU2IX1_28 ( .gnd!(gnd!), .vdd!(vdd!), .IN0(_1395_), .IN1(_1392_), .Q(_1396_), .S(_1240__bF_buf6) );
MU2X1 MU2X1_177 ( .gnd!(gnd!), .vdd!(vdd!), .IN0(_1389_), .IN1(_1396_), .Q(_1397_), .S(_1252__bF_buf3) );
AN211X1 AN211X1_2 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1226__bF_buf2), .B(_1397_), .C(_1221__bF_buf4), .D(_1382_), .Q(_1398_) );
AN311X1 AN311X1_1 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1221__bF_buf4), .B(_1364_), .C(_1367_), .D(_866__bF_buf1), .E(_1398_), .Q(_1399_) );
INX1 INX1_92 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1322__bF_buf2), .Q(_1400_) );
NO2X1 NO2X1_113 ( .gnd!(gnd!), .vdd!(vdd!), .A(_963_), .B(_1235__bF_buf0), .Q(_1401_) );
ON21X1 ON21X1_192 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1080_), .B(_1242__bF_buf3), .C(_1371_), .Q(_1402_) );
MU2IX1 MU2IX1_29 ( .gnd!(gnd!), .vdd!(vdd!), .IN0(_1402_), .IN1(_1401_), .Q(_1403_), .S(_1240__bF_buf0) );
NA2I1X1 NA2I1X1_39 ( .gnd!(gnd!), .vdd!(vdd!), .AN(_1403_), .B(_1252__bF_buf4), .Q(_1404_) );
NO3X1 NO3X1_3 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1404_), .B(_1226__bF_buf5), .C(_1400_), .Q(_1405_) );
INX1 INX1_93 ( .gnd!(gnd!), .vdd!(vdd!), .A(ALU_a_2_), .Q(_1406_) );
ON21X1 ON21X1_193 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1048__bF_buf4), .B(_931__bF_buf2), .C(ALU_b_2_), .Q(_1407_) );
NA3I1X1 NA3I1X1_8 ( .gnd!(gnd!), .vdd!(vdd!), .AN(ALU_b_2_), .B(_1143__bF_buf3), .C(_1203__bF_buf0), .Q(_1408_) );
NA3I1X1 NA3I1X1_9 ( .gnd!(gnd!), .vdd!(vdd!), .AN(_1406_), .B(_1407_), .C(_1408_), .Q(_1409_) );
INX1 INX1_94 ( .gnd!(gnd!), .vdd!(vdd!), .A(ALU_b_2_), .Q(_1410_) );
ON21X1 ON21X1_194 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1048__bF_buf4), .B(_931__bF_buf2), .C(_1410_), .Q(_1411_) );
NA3I1X1 NA3I1X1_10 ( .gnd!(gnd!), .vdd!(vdd!), .AN(_1410_), .B(_1143__bF_buf3), .C(_1203__bF_buf1), .Q(_1412_) );
NA3I1X1 NA3I1X1_11 ( .gnd!(gnd!), .vdd!(vdd!), .AN(ALU_a_2_), .B(_1411_), .C(_1412_), .Q(_1413_) );
NA2X1 NA2X1_264 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1409_), .B(_1413_), .Q(_1414_) );
AN21X1 AN21X1_81 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1208_), .B(_1207_), .C(_1080_), .Q(_1415_) );
AN21X1 AN21X1_82 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1069_), .B(_1209_), .C(_1415_), .Q(_1416_) );
NO2X1 NO2X1_114 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1414_), .B(_1416_), .Q(_1417_) );
EN3X1 EN3X1_1 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1212__bF_buf0), .B(_1406_), .C(ALU_b_2_), .Q(_1418_) );
AN21X1 AN21X1_83 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1204_), .B(_1091_), .C(ALU_a_1_), .Q(_1419_) );
ON21X1 ON21X1_195 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1419_), .B(_1213_), .C(_1205_), .Q(_1420_) );
NO2X1 NO2X1_115 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1418_), .B(_1420_), .Q(_1421_) );
ON21X1 ON21X1_196 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1421_), .B(_1417_), .C(_952__bF_buf4), .Q(_1422_) );
ON31X1 ON31X1_34 ( .gnd!(gnd!), .vdd!(vdd!), .A(_952__bF_buf5), .B(_1405_), .C(_1399_), .D(_1422_), .Q(_1423_) );
AN21X1 AN21X1_84 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1406_), .B(_1410_), .C(_1330_), .Q(_1424_) );
ON31X1 ON31X1_35 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1406_), .B(_1410_), .C(_1328__bF_buf0), .D(_1424_), .Q(_1425_) );
AN31X1 AN31X1_36 ( .gnd!(gnd!), .vdd!(vdd!), .A(ALU_a_2_), .B(ALU_b_2_), .C(_1330_), .D(_909__bF_buf0), .Q(_1426_) );
AN221X1 AN221X1_2 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1425_), .B(_1426_), .C(_1423_), .D(_909__bF_buf0), .E(_931__bF_buf3), .Q(ALU_r_2_) );
MU2IX1 MU2IX1_30 ( .gnd!(gnd!), .vdd!(vdd!), .IN0(_1254_), .IN1(_1236_), .Q(_1427_), .S(_1233__bF_buf2) );
NA2X1 NA2X1_265 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1427_), .B(_1230__bF_buf4), .Q(_1428_) );
MU2X1 MU2X1_178 ( .gnd!(gnd!), .vdd!(vdd!), .IN0(_1245_), .IN1(_1237_), .Q(_1429_), .S(_1240__bF_buf1) );
ON211X1 ON211X1_37 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1230__bF_buf3), .B(_1429_), .C(_1428_), .D(_1227__bF_buf4), .Q(_1430_) );
MU2IX1 MU2IX1_31 ( .gnd!(gnd!), .vdd!(vdd!), .IN0(_1258_), .IN1(_1253_), .Q(_1431_), .S(_1233__bF_buf2) );
NA2X1 NA2X1_266 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1431_), .B(_1252__bF_buf5), .Q(_1432_) );
NA2X1 NA2X1_267 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1230__bF_buf3), .B(ALU_a_31_), .Q(_1433_) );
NA2X1 NA2X1_268 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1432_), .B(_1433_), .Q(_1434_) );
ON21X1 ON21X1_197 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1227__bF_buf4), .B(_1434_), .C(_1430_), .Q(_1435_) );
NA2X1 NA2X1_269 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1233__bF_buf2), .B(_1266_), .Q(_1436_) );
INX1 INX1_95 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1436_), .Q(_1437_) );
MU2IX1 MU2IX1_32 ( .gnd!(gnd!), .vdd!(vdd!), .IN0(_1431_), .IN1(_1437_), .Q(_1438_), .S(_1230__bF_buf3) );
NA2X1 NA2X1_270 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1438_), .B(_1226__bF_buf4), .Q(_1439_) );
NA2X1 NA2X1_271 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1439_), .B(_1430_), .Q(_1440_) );
MU2IX1 MU2IX1_33 ( .gnd!(gnd!), .vdd!(vdd!), .IN0(_1440_), .IN1(_1435_), .Q(_1441_), .S(ALU_func7_5_bF_buf0) );
MU2IX1 MU2IX1_34 ( .gnd!(gnd!), .vdd!(vdd!), .IN0(_1249_), .IN1(_1275_), .Q(_1442_), .S(_1233__bF_buf1) );
MU2IX1 MU2IX1_35 ( .gnd!(gnd!), .vdd!(vdd!), .IN0(_1286_), .IN1(_1280_), .Q(_1443_), .S(_1240__bF_buf5) );
MU2X1 MU2X1_179 ( .gnd!(gnd!), .vdd!(vdd!), .IN0(_1442_), .IN1(_1443_), .Q(_1444_), .S(_1252__bF_buf1) );
NA2X1 NA2X1_272 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1444_), .B(_1226__bF_buf3), .Q(_1445_) );
MU2IX1 MU2IX1_36 ( .gnd!(gnd!), .vdd!(vdd!), .IN0(_1299_), .IN1(_1313_), .Q(_1446_), .S(_1240__bF_buf3) );
MU2IX1 MU2IX1_37 ( .gnd!(gnd!), .vdd!(vdd!), .IN0(_1308_), .IN1(_1291_), .Q(_1447_), .S(_1240__bF_buf3) );
MU2IX1 MU2IX1_38 ( .gnd!(gnd!), .vdd!(vdd!), .IN0(_1446_), .IN1(_1447_), .Q(_1448_), .S(_1230__bF_buf5) );
ON211X1 ON211X1_38 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1226__bF_buf2), .B(_1448_), .C(_1445_), .D(_1222__bF_buf0), .Q(_1449_) );
ON211X1 ON211X1_39 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1222__bF_buf3), .B(_1441_), .C(_1449_), .D(EXT_type_bF_buf1), .Q(_1450_) );
NA2I1X1 NA2I1X1_40 ( .gnd!(gnd!), .vdd!(vdd!), .AN(_1300_), .B(_1296_), .Q(_1451_) );
MU2IX1 MU2IX1_39 ( .gnd!(gnd!), .vdd!(vdd!), .IN0(_1451_), .IN1(_1318_), .Q(_1452_), .S(_1240__bF_buf0) );
NA2X1 NA2X1_273 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1452_), .B(_1252__bF_buf4), .Q(_1453_) );
NA2I1X1 NA2I1X1_41 ( .gnd!(gnd!), .vdd!(vdd!), .AN(_1453_), .B(_1227__bF_buf5), .Q(_1454_) );
NO2X1 NO2X1_116 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1400_), .B(_1454_), .Q(_1455_) );
NO2X1 NO2X1_117 ( .gnd!(gnd!), .vdd!(vdd!), .A(_952__bF_buf5), .B(_1455_), .Q(_1456_) );
INX1 INX1_96 ( .gnd!(gnd!), .vdd!(vdd!), .A(ALU_b_3_), .Q(_1457_) );
ON21X1 ON21X1_198 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1048__bF_buf1), .B(_931__bF_buf4), .C(_1457_), .Q(_1458_) );
NA3I1X1 NA3I1X1_12 ( .gnd!(gnd!), .vdd!(vdd!), .AN(_1457_), .B(_1143__bF_buf3), .C(_1203__bF_buf1), .Q(_1459_) );
AN21X1 AN21X1_85 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1459_), .B(_1458_), .C(_1295_), .Q(_1460_) );
ON21X1 ON21X1_199 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1048__bF_buf1), .B(_931__bF_buf4), .C(ALU_b_3_), .Q(_1461_) );
NA3I1X1 NA3I1X1_13 ( .gnd!(gnd!), .vdd!(vdd!), .AN(ALU_b_3_), .B(_1143__bF_buf3), .C(_1203__bF_buf1), .Q(_1462_) );
AN21X1 AN21X1_86 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1462_), .B(_1461_), .C(ALU_a_3_), .Q(_1463_) );
ON221X1 ON221X1_1 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1460_), .B(_1463_), .C(_1414_), .D(_1416_), .E(_1409_), .Q(_1464_) );
EN3X1 EN3X1_2 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1212__bF_buf0), .B(_1295_), .C(ALU_b_3_), .Q(_1465_) );
ON21X1 ON21X1_200 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1416_), .B(_1414_), .C(_1409_), .Q(_1466_) );
NA2X1 NA2X1_274 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1466_), .B(_1465_), .Q(_1467_) );
NA2X1 NA2X1_275 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1467_), .B(_1464_), .Q(_1468_) );
AO22X2 AO22X2_23 ( .gnd!(gnd!), .vdd!(vdd!), .A(_952__bF_buf1), .B(_1468_), .C(_1450_), .D(_1456_), .Q(_1469_) );
AN21X1 AN21X1_87 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1295_), .B(_1457_), .C(_1330_), .Q(_1470_) );
ON31X1 ON31X1_36 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1295_), .B(_1457_), .C(_1328__bF_buf0), .D(_1470_), .Q(_1471_) );
AN31X1 AN31X1_37 ( .gnd!(gnd!), .vdd!(vdd!), .A(ALU_a_3_), .B(ALU_b_3_), .C(_1330_), .D(_909__bF_buf2), .Q(_1472_) );
AN221X1 AN221X1_3 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1471_), .B(_1472_), .C(_1469_), .D(_909__bF_buf2), .E(_931__bF_buf3), .Q(ALU_r_3_) );
INX1 INX1_97 ( .gnd!(gnd!), .vdd!(vdd!), .A(ALU_b_4_), .Q(_1473_) );
ON21X1 ON21X1_201 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1048__bF_buf4), .B(_931__bF_buf2), .C(_1473_), .Q(_1474_) );
NA3I1X1 NA3I1X1_14 ( .gnd!(gnd!), .vdd!(vdd!), .AN(_1473_), .B(_1143__bF_buf3), .C(_1203__bF_buf1), .Q(_1475_) );
AN21X1 AN21X1_88 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1475_), .B(_1474_), .C(_1297_), .Q(_1476_) );
ON21X1 ON21X1_202 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1048__bF_buf3), .B(_931__bF_buf1), .C(ALU_b_4_), .Q(_1477_) );
NA3I1X1 NA3I1X1_15 ( .gnd!(gnd!), .vdd!(vdd!), .AN(ALU_b_4_), .B(_1143__bF_buf2), .C(_1203__bF_buf0), .Q(_1478_) );
AN21X1 AN21X1_89 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1478_), .B(_1477_), .C(ALU_a_4_), .Q(_1479_) );
NO2X1 NO2X1_118 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1476_), .B(_1479_), .Q(_1480_) );
NA2X1 NA2X1_276 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1412_), .B(_1411_), .Q(_1481_) );
NA3I1X1 NA3I1X1_16 ( .gnd!(gnd!), .vdd!(vdd!), .AN(ALU_a_3_), .B(_1458_), .C(_1459_), .Q(_1482_) );
AN31X1 AN31X1_38 ( .gnd!(gnd!), .vdd!(vdd!), .A(ALU_a_2_), .B(_1481_), .C(_1482_), .D(_1460_), .Q(_1483_) );
AN21X1 AN21X1_90 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1459_), .B(_1458_), .C(ALU_a_3_), .Q(_1484_) );
AN21X1 AN21X1_91 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1462_), .B(_1461_), .C(_1295_), .Q(_1485_) );
ON211X1 ON211X1_40 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1484_), .B(_1485_), .C(_1409_), .D(_1413_), .Q(_1486_) );
ON21X1 ON21X1_203 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1486_), .B(_1416_), .C(_1483_), .Q(_1487_) );
NA2X1 NA2X1_277 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1487_), .B(_1480_), .Q(_1488_) );
NA3I1X1 NA3I1X1_17 ( .gnd!(gnd!), .vdd!(vdd!), .AN(_1295_), .B(_1461_), .C(_1462_), .Q(_1489_) );
ON21X1 ON21X1_204 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1463_), .B(_1409_), .C(_1489_), .Q(_1490_) );
AN31X1 AN31X1_39 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1418_), .B(_1465_), .C(_1420_), .D(_1490_), .Q(_1491_) );
NA2I1X1 NA2I1X1_42 ( .gnd!(gnd!), .vdd!(vdd!), .AN(_1480_), .B(_1491_), .Q(_1492_) );
NA2X1 NA2X1_278 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1492_), .B(_1488_), .Q(_1493_) );
NA2X1 NA2X1_279 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1493_), .B(_952__bF_buf4), .Q(_1494_) );
NA2X1 NA2X1_280 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1433_), .B(_1226__bF_buf4), .Q(_1495_) );
MU2IX1 MU2IX1_40 ( .gnd!(gnd!), .vdd!(vdd!), .IN0(_1336_), .IN1(_1355_), .Q(_1496_), .S(_1240__bF_buf5) );
MU2IX1 MU2IX1_41 ( .gnd!(gnd!), .vdd!(vdd!), .IN0(_1343_), .IN1(_1339_), .Q(_1497_), .S(_1240__bF_buf5) );
MU2IX1 MU2IX1_42 ( .gnd!(gnd!), .vdd!(vdd!), .IN0(_1496_), .IN1(_1497_), .Q(_1498_), .S(_1252__bF_buf3) );
MU2IX1 MU2IX1_43 ( .gnd!(gnd!), .vdd!(vdd!), .IN0(_1351_), .IN1(_1360_), .Q(_1499_), .S(_1240__bF_buf1) );
NO2X1 NO2X1_119 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1230__bF_buf5), .B(_1499_), .Q(_1500_) );
ON22X1 ON22X1_2 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1498_), .B(_1226__bF_buf3), .C(_1500_), .D(_1495_), .Q(_1501_) );
MU2IX1 MU2IX1_44 ( .gnd!(gnd!), .vdd!(vdd!), .IN0(_1498_), .IN1(_1500_), .Q(_1502_), .S(_1226__bF_buf3) );
MU2IX1 MU2IX1_45 ( .gnd!(gnd!), .vdd!(vdd!), .IN0(_1502_), .IN1(_1501_), .Q(_1503_), .S(ALU_func7_5_bF_buf0) );
NO2X1 NO2X1_120 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1222__bF_buf0), .B(_1503_), .Q(_1504_) );
MU2IX1 MU2IX1_46 ( .gnd!(gnd!), .vdd!(vdd!), .IN0(_1385_), .IN1(_1346_), .Q(_1505_), .S(_1240__bF_buf4) );
MU2X1 MU2X1_180 ( .gnd!(gnd!), .vdd!(vdd!), .IN0(_1388_), .IN1(_1392_), .Q(_1506_), .S(_1233__bF_buf4) );
MU2IX1 MU2IX1_47 ( .gnd!(gnd!), .vdd!(vdd!), .IN0(_1506_), .IN1(_1505_), .Q(_1507_), .S(_1230__bF_buf1) );
MU2X1 MU2X1_181 ( .gnd!(gnd!), .vdd!(vdd!), .IN0(_1395_), .IN1(_1376_), .Q(_1508_), .S(_1233__bF_buf4) );
NA2X1 NA2X1_281 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1379_), .B(_1240__bF_buf6), .Q(_1509_) );
ON21X1 ON21X1_205 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1370_), .B(_1240__bF_buf6), .C(_1509_), .Q(_1510_) );
MU2IX1 MU2IX1_48 ( .gnd!(gnd!), .vdd!(vdd!), .IN0(_1510_), .IN1(_1508_), .Q(_1511_), .S(_1230__bF_buf1) );
MU2IX1 MU2IX1_49 ( .gnd!(gnd!), .vdd!(vdd!), .IN0(_1507_), .IN1(_1511_), .Q(_1512_), .S(_1227__bF_buf6) );
AN211X1 AN211X1_3 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1222__bF_buf3), .B(_1512_), .C(_866__bF_buf4), .D(_1504_), .Q(_1513_) );
AND2X2 AND2X2_6 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1233__bF_buf0), .B(_1401_), .Q(_1514_) );
MU2IX1 MU2IX1_50 ( .gnd!(gnd!), .vdd!(vdd!), .IN0(_1297_), .IN1(_1295_), .Q(_1515_), .S(_1235__bF_buf0) );
MU2X1 MU2X1_182 ( .gnd!(gnd!), .vdd!(vdd!), .IN0(_1515_), .IN1(_1402_), .Q(_1516_), .S(_1240__bF_buf0) );
MU2IX1 MU2IX1_51 ( .gnd!(gnd!), .vdd!(vdd!), .IN0(_1516_), .IN1(_1514_), .Q(_1517_), .S(_1230__bF_buf2) );
NO2X1 NO2X1_121 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1226__bF_buf5), .B(_1517_), .Q(_1518_) );
AND2X2 AND2X2_7 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1518_), .B(_1322__bF_buf2), .Q(_1519_) );
ON31X1 ON31X1_37 ( .gnd!(gnd!), .vdd!(vdd!), .A(_952__bF_buf1), .B(_1519_), .C(_1513_), .D(_1494_), .Q(_1520_) );
AN21X1 AN21X1_92 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1297_), .B(_1473_), .C(_1330_), .Q(_1521_) );
ON31X1 ON31X1_38 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1297_), .B(_1473_), .C(_1328__bF_buf4), .D(_1521_), .Q(_1522_) );
AN31X1 AN31X1_40 ( .gnd!(gnd!), .vdd!(vdd!), .A(ALU_a_4_), .B(ALU_b_4_), .C(_1330_), .D(_909__bF_buf0), .Q(_1523_) );
AN221X1 AN221X1_4 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1522_), .B(_1523_), .C(_1520_), .D(_909__bF_buf0), .E(_931__bF_buf3), .Q(ALU_r_4_) );
NO2X2 NO2X2_2 ( .gnd!(gnd!), .vdd!(vdd!), .A(_920_), .B(_888__bF_buf4), .Q(_1524_) );
INX2 INX2_9 ( .gnd!(gnd!), .vdd!(vdd!), .A(_909__bF_buf1), .Q(_1525_) );
INX2 INX2_10 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1330_), .Q(_1526_) );
NA2X1 NA2X1_282 ( .gnd!(gnd!), .vdd!(vdd!), .A(ALU_a_5_), .B(ALU_b_5_), .Q(_1527_) );
NO2X1 NO2X1_122 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1527_), .B(_1328__bF_buf3), .Q(_1528_) );
ON22X1 ON22X1_3 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1329__bF_buf4), .B(_888__bF_buf1), .C(ALU_a_5_), .D(ALU_b_5_), .Q(_1529_) );
ON22X1 ON22X1_4 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1528_), .B(_1529_), .C(_1526__bF_buf1), .D(_1527_), .Q(_1530_) );
NA2X1 NA2X1_283 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1530_), .B(_1525__bF_buf3), .Q(_1531_) );
NA2X1 NA2X1_284 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1255_), .B(_1230__bF_buf4), .Q(_1532_) );
NA2X1 NA2X1_285 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1238_), .B(_1252__bF_buf5), .Q(_1533_) );
AND3X4 AND3X4_1 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1532_), .B(_1533_), .C(_1227__bF_buf2), .Q(_1534_) );
NO2X1 NO2X1_123 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1230__bF_buf4), .B(_1267_), .Q(_1535_) );
NO2X1 NO2X1_124 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1227__bF_buf2), .B(_1535_), .Q(_1536_) );
NO3X1 NO3X1_4 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1534_), .B(ALU_func7_5_bF_buf2), .C(_1536_), .Q(_1537_) );
NA2X1 NA2X1_286 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1260_), .B(_1252__bF_buf5), .Q(_1538_) );
AN31X1 AN31X1_41 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1226__bF_buf1), .B(_1433_), .C(_1538_), .D(_1534_), .Q(_1539_) );
AND2X2 AND2X2_8 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1539_), .B(ALU_func7_5_bF_buf2), .Q(_1540_) );
MU2X1 MU2X1_183 ( .gnd!(gnd!), .vdd!(vdd!), .IN0(_1314_), .IN1(_1292_), .Q(_1541_), .S(_1230__bF_buf3) );
NA2X1 NA2X1_287 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1541_), .B(_1227__bF_buf2), .Q(_1542_) );
NA2X1 NA2X1_288 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1250_), .B(_1230__bF_buf4), .Q(_1543_) );
ON21X1 ON21X1_206 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1281_), .B(_1230__bF_buf4), .C(_1543_), .Q(_1544_) );
ON211X1 ON211X1_41 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1544_), .B(_1227__bF_buf2), .C(_1222__bF_buf5), .D(_1542_), .Q(_1545_) );
ON311X1 ON311X1_1 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1222__bF_buf5), .B(_1537_), .C(_1540_), .D(EXT_type_bF_buf4), .E(_1545_), .Q(_1546_) );
NA2X1 NA2X1_289 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1310_), .B(_1298_), .Q(_1547_) );
MU2IX1 MU2IX1_52 ( .gnd!(gnd!), .vdd!(vdd!), .IN0(_1451_), .IN1(_1547_), .Q(_1548_), .S(_1233__bF_buf0) );
MU2IX1 MU2IX1_53 ( .gnd!(gnd!), .vdd!(vdd!), .IN0(_1548_), .IN1(_1319_), .Q(_1549_), .S(_1230__bF_buf2) );
NO2X1 NO2X1_125 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1226__bF_buf5), .B(_1549_), .Q(_1550_) );
NA2X1 NA2X1_290 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1550_), .B(_1322__bF_buf2), .Q(_1551_) );
INX1 INX1_98 ( .gnd!(gnd!), .vdd!(vdd!), .A(ALU_b_5_), .Q(_1552_) );
ON21X1 ON21X1_207 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1048__bF_buf3), .B(_931__bF_buf1), .C(_1552_), .Q(_1553_) );
NA3I1X1 NA3I1X1_18 ( .gnd!(gnd!), .vdd!(vdd!), .AN(_1552_), .B(_1143__bF_buf2), .C(_1203__bF_buf0), .Q(_1554_) );
AN21X1 AN21X1_93 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1554_), .B(_1553_), .C(_1309_), .Q(_1555_) );
ON21X1 ON21X1_208 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1048__bF_buf4), .B(_931__bF_buf2), .C(ALU_b_5_), .Q(_1556_) );
NA3I1X1 NA3I1X1_19 ( .gnd!(gnd!), .vdd!(vdd!), .AN(ALU_b_5_), .B(_1143__bF_buf2), .C(_1203__bF_buf0), .Q(_1557_) );
AN21X1 AN21X1_94 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1557_), .B(_1556_), .C(ALU_a_5_), .Q(_1558_) );
NO2X1 NO2X1_126 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1555_), .B(_1558_), .Q(_1559_) );
AN211X1 AN211X1_4 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1480_), .B(_1487_), .C(_1476_), .D(_1559_), .Q(_1560_) );
NA3I1X1 NA3I1X1_20 ( .gnd!(gnd!), .vdd!(vdd!), .AN(_1297_), .B(_1477_), .C(_1478_), .Q(_1561_) );
INX1 INX1_99 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1559_), .Q(_1562_) );
AN21X1 AN21X1_95 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1488_), .B(_1561_), .C(_1562_), .Q(_1563_) );
NO2X1 NO2X1_127 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1560_), .B(_1563_), .Q(_1564_) );
NO2X1 NO2X1_128 ( .gnd!(gnd!), .vdd!(vdd!), .A(_941__bF_buf2), .B(_1564_), .Q(_1565_) );
AO311X1 AO311X1_1 ( .gnd!(gnd!), .vdd!(vdd!), .A(_941__bF_buf3), .B(_1551_), .C(_1546_), .D(_1525__bF_buf2), .E(_1565_), .Q(_1566_) );
AN22X1 AN22X1_22 ( .gnd!(gnd!), .vdd!(vdd!), .A(_866__bF_buf0), .B(_1524__bF_buf0), .C(_1566_), .D(_1531_), .Q(ALU_r_5_) );
NA2X1 NA2X1_291 ( .gnd!(gnd!), .vdd!(vdd!), .A(ALU_a_6_), .B(ALU_b_6_), .Q(_1567_) );
NO2X1 NO2X1_129 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1567_), .B(_1328__bF_buf3), .Q(_1568_) );
ON22X1 ON22X1_5 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1329__bF_buf4), .B(_888__bF_buf1), .C(ALU_a_6_), .D(ALU_b_6_), .Q(_1569_) );
ON22X1 ON22X1_6 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1568_), .B(_1569_), .C(_1526__bF_buf0), .D(_1567_), .Q(_1570_) );
NA2X1 NA2X1_292 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1570_), .B(_1525__bF_buf3), .Q(_1571_) );
NA2X1 NA2X1_293 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1357_), .B(_1230__bF_buf5), .Q(_1572_) );
NA2X1 NA2X1_294 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1340_), .B(_1252__bF_buf1), .Q(_1573_) );
AND3X4 AND3X4_2 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1573_), .B(_1227__bF_buf6), .C(_1572_), .Q(_1574_) );
AND2X2 AND2X2_9 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1259_), .B(_1433_), .Q(_1575_) );
NO2X1 NO2X1_130 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1575_), .B(_1574_), .Q(_1576_) );
AND2X2 AND2X2_10 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1576_), .B(ALU_func7_5_bF_buf1), .Q(_1577_) );
NA2I1X1 NA2I1X1_43 ( .gnd!(gnd!), .vdd!(vdd!), .AN(_1361_), .B(_1252__bF_buf5), .Q(_1578_) );
AN21X1 AN21X1_96 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1226__bF_buf2), .B(_1578_), .C(_1574_), .Q(_1579_) );
MU2X1 MU2X1_184 ( .gnd!(gnd!), .vdd!(vdd!), .IN0(_1396_), .IN1(_1380_), .Q(_1580_), .S(_1252__bF_buf3) );
NA2X1 NA2X1_295 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1580_), .B(_1227__bF_buf6), .Q(_1581_) );
MU2IX1 MU2IX1_54 ( .gnd!(gnd!), .vdd!(vdd!), .IN0(_1347_), .IN1(_1389_), .Q(_1582_), .S(_1252__bF_buf1) );
ON211X1 ON211X1_42 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1227__bF_buf6), .B(_1582_), .C(_1581_), .D(_1222__bF_buf0), .Q(_1583_) );
ON311X1 ON311X1_2 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1222__bF_buf2), .B(_1579_), .C(_1577_), .D(EXT_type_bF_buf1), .E(_1583_), .Q(_1584_) );
AND2X2 AND2X2_11 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1377_), .B(_1369_), .Q(_1585_) );
MU2IX1 MU2IX1_55 ( .gnd!(gnd!), .vdd!(vdd!), .IN0(_1585_), .IN1(_1515_), .Q(_1586_), .S(_1240__bF_buf0) );
MU2X1 MU2X1_185 ( .gnd!(gnd!), .vdd!(vdd!), .IN0(_1586_), .IN1(_1403_), .Q(_1587_), .S(_1230__bF_buf2) );
ON31X1 ON31X1_39 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1226__bF_buf5), .B(_1400_), .C(_1587_), .D(_1584_), .Q(_1588_) );
NA3I1X1 NA3I1X1_21 ( .gnd!(gnd!), .vdd!(vdd!), .AN(ALU_a_5_), .B(_1553_), .C(_1554_), .Q(_1589_) );
ON21X1 ON21X1_209 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1476_), .B(_1555_), .C(_1589_), .Q(_1590_) );
NA3I1X1 NA3I1X1_22 ( .gnd!(gnd!), .vdd!(vdd!), .AN(ALU_a_4_), .B(_1474_), .C(_1475_), .Q(_1591_) );
AN21X1 AN21X1_97 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1554_), .B(_1553_), .C(ALU_a_5_), .Q(_1592_) );
AN21X1 AN21X1_98 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1557_), .B(_1556_), .C(_1309_), .Q(_1593_) );
ON211X1 ON211X1_43 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1592_), .B(_1593_), .C(_1561_), .D(_1591_), .Q(_1594_) );
NA2I1X1 NA2I1X1_44 ( .gnd!(gnd!), .vdd!(vdd!), .AN(_1594_), .B(_1487_), .Q(_1595_) );
ON21X1 ON21X1_210 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1048__bF_buf2), .B(_931__bF_buf5), .C(ALU_b_6_), .Q(_1596_) );
NA3I1X1 NA3I1X1_23 ( .gnd!(gnd!), .vdd!(vdd!), .AN(ALU_b_6_), .B(_1143__bF_buf0), .C(_1203__bF_buf3), .Q(_1597_) );
NA3I1X1 NA3I1X1_24 ( .gnd!(gnd!), .vdd!(vdd!), .AN(ALU_a_6_), .B(_1596_), .C(_1597_), .Q(_1598_) );
INX1 INX1_100 ( .gnd!(gnd!), .vdd!(vdd!), .A(ALU_b_6_), .Q(_1599_) );
ON21X1 ON21X1_211 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1048__bF_buf2), .B(_931__bF_buf5), .C(_1599_), .Q(_1600_) );
NA3I1X1 NA3I1X1_25 ( .gnd!(gnd!), .vdd!(vdd!), .AN(_1599_), .B(_1143__bF_buf4), .C(_1203__bF_buf3), .Q(_1601_) );
NA3I1X1 NA3I1X1_26 ( .gnd!(gnd!), .vdd!(vdd!), .AN(_1311_), .B(_1600_), .C(_1601_), .Q(_1602_) );
AN22X1 AN22X1_23 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1598_), .B(_1602_), .C(_1595_), .D(_1590_), .Q(_1603_) );
AN21X1 AN21X1_99 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1601_), .B(_1600_), .C(ALU_a_6_), .Q(_1604_) );
AN21X1 AN21X1_100 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1597_), .B(_1596_), .C(_1311_), .Q(_1605_) );
NO2X1 NO2X1_131 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1604_), .B(_1605_), .Q(_1606_) );
OA211X4 OA211X4_1 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1491_), .B(_1594_), .C(_1590_), .D(_1606_), .Q(_1607_) );
ON21X1 ON21X1_212 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1603_), .B(_1607_), .C(_952__bF_buf4), .Q(_1608_) );
ON211X1 ON211X1_44 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1588_), .B(_952__bF_buf1), .C(_909__bF_buf4), .D(_1608_), .Q(_1609_) );
AN22X1 AN22X1_24 ( .gnd!(gnd!), .vdd!(vdd!), .A(_866__bF_buf2), .B(_1524__bF_buf3), .C(_1609_), .D(_1571_), .Q(ALU_r_6_) );
NA2X1 NA2X1_296 ( .gnd!(gnd!), .vdd!(vdd!), .A(ALU_a_7_), .B(ALU_b_7_), .Q(_1610_) );
NO2X1 NO2X1_132 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1610_), .B(_1328__bF_buf4), .Q(_1611_) );
ON22X1 ON22X1_7 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1329__bF_buf4), .B(_888__bF_buf2), .C(ALU_a_7_), .D(ALU_b_7_), .Q(_1612_) );
ON22X1 ON22X1_8 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1611_), .B(_1612_), .C(_1526__bF_buf2), .D(_1610_), .Q(_1613_) );
NA2X1 NA2X1_297 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1613_), .B(_1525__bF_buf4), .Q(_1614_) );
NA3I1X1 NA3I1X1_27 ( .gnd!(gnd!), .vdd!(vdd!), .AN(_1309_), .B(_1556_), .C(_1557_), .Q(_1615_) );
AN21X1 AN21X1_101 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1561_), .B(_1615_), .C(_1558_), .Q(_1616_) );
AN31X1 AN31X1_42 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1480_), .B(_1559_), .C(_1487_), .D(_1616_), .Q(_1617_) );
NA3I1X1 NA3I1X1_28 ( .gnd!(gnd!), .vdd!(vdd!), .AN(_1311_), .B(_1596_), .C(_1597_), .Q(_1618_) );
ON21X1 ON21X1_213 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1048__bF_buf3), .B(_931__bF_buf1), .C(ALU_b_7_), .Q(_1619_) );
NA3I1X1 NA3I1X1_29 ( .gnd!(gnd!), .vdd!(vdd!), .AN(ALU_b_7_), .B(_1143__bF_buf0), .C(_1203__bF_buf3), .Q(_1620_) );
NA3I1X1 NA3I1X1_30 ( .gnd!(gnd!), .vdd!(vdd!), .AN(ALU_a_7_), .B(_1619_), .C(_1620_), .Q(_1621_) );
INX1 INX1_101 ( .gnd!(gnd!), .vdd!(vdd!), .A(ALU_b_7_), .Q(_1622_) );
ON21X1 ON21X1_214 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1048__bF_buf2), .B(_931__bF_buf5), .C(_1622_), .Q(_1623_) );
NA3I1X1 NA3I1X1_31 ( .gnd!(gnd!), .vdd!(vdd!), .AN(_1622_), .B(_1143__bF_buf0), .C(_1203__bF_buf3), .Q(_1624_) );
NA3I1X1 NA3I1X1_32 ( .gnd!(gnd!), .vdd!(vdd!), .AN(_1304_), .B(_1623_), .C(_1624_), .Q(_1625_) );
NA2X1 NA2X1_298 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1621_), .B(_1625_), .Q(_1626_) );
INX1 INX1_102 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1626_), .Q(_1627_) );
ON211X1 ON211X1_45 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1617_), .B(_1606_), .C(_1627_), .D(_1618_), .Q(_1628_) );
ON21X1 ON21X1_215 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1617_), .B(_1606_), .C(_1618_), .Q(_1629_) );
NA2X1 NA2X1_299 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1629_), .B(_1626_), .Q(_1630_) );
NA2X1 NA2X1_300 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1630_), .B(_1628_), .Q(_1631_) );
NA2X1 NA2X1_301 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1631_), .B(_952__bF_buf4), .Q(_1632_) );
NA2X1 NA2X1_302 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1431_), .B(_1230__bF_buf3), .Q(_1633_) );
NA2X1 NA2X1_303 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1427_), .B(_1252__bF_buf5), .Q(_1634_) );
NA2X1 NA2X1_304 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1633_), .B(_1634_), .Q(_1635_) );
NO2X1 NO2X1_133 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1226__bF_buf4), .B(_1635_), .Q(_1636_) );
NO2X1 NO2X1_134 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1230__bF_buf5), .B(_1436_), .Q(_1637_) );
NO2X1 NO2X1_135 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1227__bF_buf1), .B(_1637_), .Q(_1638_) );
NO2X1 NO2X1_136 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1638_), .B(_1636_), .Q(_1639_) );
NA2X1 NA2X1_305 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1639_), .B(_1223_), .Q(_1640_) );
NO2X1 NO2X1_137 ( .gnd!(gnd!), .vdd!(vdd!), .A(ALU_a_31_), .B(_1227__bF_buf1), .Q(_1641_) );
OR2X2 OR2X2_12 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1636_), .B(_1641_), .Q(_1642_) );
NA2I1X1 NA2I1X1_45 ( .gnd!(gnd!), .vdd!(vdd!), .AN(_1642_), .B(ALU_func7_5_bF_buf1), .Q(_1643_) );
MU2IX1 MU2IX1_56 ( .gnd!(gnd!), .vdd!(vdd!), .IN0(_1443_), .IN1(_1447_), .Q(_1644_), .S(_1252__bF_buf1) );
NA2X1 NA2X1_306 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1442_), .B(_1252__bF_buf1), .Q(_1645_) );
ON21X1 ON21X1_216 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1252__bF_buf1), .B(_1429_), .C(_1645_), .Q(_1646_) );
NA2X1 NA2X1_307 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1646_), .B(_1226__bF_buf3), .Q(_1647_) );
OA211X4 OA211X4_2 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1226__bF_buf3), .B(_1644_), .C(_1647_), .D(_1222__bF_buf0), .Q(_1648_) );
AN311X1 AN311X1_2 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1221__bF_buf4), .B(_1640_), .C(_1643_), .D(_866__bF_buf1), .E(_1648_), .Q(_1649_) );
NA2X1 NA2X1_308 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1305_), .B(_1312_), .Q(_1650_) );
MU2IX1 MU2IX1_57 ( .gnd!(gnd!), .vdd!(vdd!), .IN0(_1650_), .IN1(_1547_), .Q(_1651_), .S(_1240__bF_buf6) );
MU2X1 MU2X1_186 ( .gnd!(gnd!), .vdd!(vdd!), .IN0(_1452_), .IN1(_1651_), .Q(_1652_), .S(_1252__bF_buf4) );
NA2X1 NA2X1_309 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1652_), .B(_1227__bF_buf5), .Q(_1653_) );
NO2X1 NO2X1_138 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1400_), .B(_1653_), .Q(_1654_) );
ON311X1 ON311X1_3 ( .gnd!(gnd!), .vdd!(vdd!), .A(_952__bF_buf5), .B(_1654_), .C(_1649_), .D(_909__bF_buf3), .E(_1632_), .Q(_1655_) );
AN22X1 AN22X1_25 ( .gnd!(gnd!), .vdd!(vdd!), .A(_866__bF_buf0), .B(_1524__bF_buf0), .C(_1655_), .D(_1614_), .Q(ALU_r_7_) );
NA2X1 NA2X1_310 ( .gnd!(gnd!), .vdd!(vdd!), .A(ALU_a_8_), .B(ALU_b_8_), .Q(_1656_) );
NO2X1 NO2X1_139 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1656_), .B(_1328__bF_buf3), .Q(_1657_) );
ON22X1 ON22X1_9 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1329__bF_buf4), .B(_888__bF_buf1), .C(ALU_a_8_), .D(ALU_b_8_), .Q(_1658_) );
ON22X1 ON22X1_10 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1657_), .B(_1658_), .C(_1526__bF_buf2), .D(_1656_), .Q(_1659_) );
NA2X1 NA2X1_311 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1659_), .B(_1525__bF_buf0), .Q(_1660_) );
ON21X1 ON21X1_217 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1048__bF_buf1), .B(_931__bF_buf4), .C(ALU_b_8_), .Q(_1661_) );
NA3I1X1 NA3I1X1_33 ( .gnd!(gnd!), .vdd!(vdd!), .AN(ALU_b_8_), .B(_1143__bF_buf2), .C(_1203__bF_buf4), .Q(_1662_) );
NA3I1X1 NA3I1X1_34 ( .gnd!(gnd!), .vdd!(vdd!), .AN(_1306_), .B(_1661_), .C(_1662_), .Q(_1663_) );
INX1 INX1_103 ( .gnd!(gnd!), .vdd!(vdd!), .A(ALU_b_8_), .Q(_1664_) );
ON21X1 ON21X1_218 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1048__bF_buf1), .B(_931__bF_buf4), .C(_1664_), .Q(_1665_) );
NA3I1X1 NA3I1X1_35 ( .gnd!(gnd!), .vdd!(vdd!), .AN(_1664_), .B(_1143__bF_buf2), .C(_1203__bF_buf4), .Q(_1666_) );
NA3I1X1 NA3I1X1_36 ( .gnd!(gnd!), .vdd!(vdd!), .AN(ALU_a_8_), .B(_1665_), .C(_1666_), .Q(_1667_) );
NA2X1 NA2X1_312 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1663_), .B(_1667_), .Q(_1668_) );
NA3I1X1 NA3I1X1_37 ( .gnd!(gnd!), .vdd!(vdd!), .AN(_1304_), .B(_1619_), .C(_1620_), .Q(_1669_) );
NA3I1X1 NA3I1X1_38 ( .gnd!(gnd!), .vdd!(vdd!), .AN(ALU_a_7_), .B(_1623_), .C(_1624_), .Q(_1670_) );
ON211X1 ON211X1_46 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1604_), .B(_1605_), .C(_1669_), .D(_1670_), .Q(_1671_) );
NO2X1 NO2X1_140 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1594_), .B(_1671_), .Q(_1672_) );
NA2X1 NA2X1_313 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1669_), .B(_1618_), .Q(_1673_) );
NA2X1 NA2X1_314 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1673_), .B(_1670_), .Q(_1674_) );
ON21X1 ON21X1_219 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1671_), .B(_1590_), .C(_1674_), .Q(_1675_) );
AN21X1 AN21X1_102 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1487_), .B(_1672_), .C(_1675_), .Q(_1676_) );
NO2X1 NO2X1_141 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1668_), .B(_1676_), .Q(_1677_) );
AN22X1 AN22X1_26 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1598_), .B(_1602_), .C(_1621_), .D(_1625_), .Q(_1678_) );
NA3X1 NA3X1_3 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1559_), .B(_1480_), .C(_1678_), .Q(_1679_) );
AN22X1 AN22X1_27 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1670_), .B(_1673_), .C(_1678_), .D(_1616_), .Q(_1680_) );
ON21X1 ON21X1_220 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1491_), .B(_1679_), .C(_1680_), .Q(_1681_) );
NO2I1X1 NO2I1X1_34 ( .gnd!(gnd!), .vdd!(vdd!), .AN(_1668_), .B(_1681_), .Q(_1682_) );
NO2X1 NO2X1_142 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1682_), .B(_1677_), .Q(_1683_) );
NA2X1 NA2X1_315 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1514_), .B(_1252__bF_buf2), .Q(_1684_) );
AND2X2 AND2X2_12 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1374_), .B(_1378_), .Q(_1685_) );
MU2X1 MU2X1_187 ( .gnd!(gnd!), .vdd!(vdd!), .IN0(_1685_), .IN1(_1585_), .Q(_1686_), .S(_1240__bF_buf6) );
MU2IX1 MU2IX1_58 ( .gnd!(gnd!), .vdd!(vdd!), .IN0(_1686_), .IN1(_1516_), .Q(_1687_), .S(_1230__bF_buf2) );
MU2IX1 MU2IX1_59 ( .gnd!(gnd!), .vdd!(vdd!), .IN0(_1687_), .IN1(_1684_), .Q(_1688_), .S(_1226__bF_buf6) );
MU2X1 MU2X1_188 ( .gnd!(gnd!), .vdd!(vdd!), .IN0(_1506_), .IN1(_1508_), .Q(_1689_), .S(_1252__bF_buf0) );
MU2IX1 MU2IX1_60 ( .gnd!(gnd!), .vdd!(vdd!), .IN0(_1497_), .IN1(_1505_), .Q(_1690_), .S(_1252__bF_buf3) );
NA2X1 NA2X1_316 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1690_), .B(_1226__bF_buf2), .Q(_1691_) );
ON211X1 ON211X1_47 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1689_), .B(_1226__bF_buf2), .C(_1222__bF_buf0), .D(_1691_), .Q(_1692_) );
MU2IX1 MU2IX1_61 ( .gnd!(gnd!), .vdd!(vdd!), .IN0(_1499_), .IN1(_1496_), .Q(_1693_), .S(_1252__bF_buf1) );
NA2X1 NA2X1_317 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1693_), .B(_1227__bF_buf6), .Q(_1694_) );
NA2X1 NA2X1_318 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1226__bF_buf1), .B(ALU_a_31_), .Q(_1695_) );
ON211X1 ON211X1_48 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1223_), .B(_1695_), .C(_1694_), .D(_1221__bF_buf4), .Q(_1696_) );
AN32X1 AN32X1_1 ( .gnd!(gnd!), .vdd!(vdd!), .A(EXT_type_bF_buf6), .B(_1696_), .C(_1692_), .D(_1322__bF_buf0), .E(_1688_), .Q(_1697_) );
NA2X1 NA2X1_319 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1697_), .B(_941__bF_buf4), .Q(_1698_) );
ON211X1 ON211X1_49 ( .gnd!(gnd!), .vdd!(vdd!), .A(_941__bF_buf0), .B(_1683_), .C(_1698_), .D(_909__bF_buf1), .Q(_1699_) );
AN22X1 AN22X1_28 ( .gnd!(gnd!), .vdd!(vdd!), .A(_866__bF_buf5), .B(_1524__bF_buf1), .C(_1699_), .D(_1660_), .Q(ALU_r_8_) );
NA2X1 NA2X1_320 ( .gnd!(gnd!), .vdd!(vdd!), .A(ALU_a_9_), .B(ALU_b_9_), .Q(_1700_) );
NO2X1 NO2X1_143 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1700_), .B(_1328__bF_buf3), .Q(_1701_) );
ON22X1 ON22X1_11 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1329__bF_buf4), .B(_888__bF_buf1), .C(ALU_a_9_), .D(ALU_b_9_), .Q(_1702_) );
ON22X1 ON22X1_12 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1701_), .B(_1702_), .C(_1526__bF_buf0), .D(_1700_), .Q(_1703_) );
NA2X1 NA2X1_321 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1703_), .B(_1525__bF_buf4), .Q(_1704_) );
NA2X1 NA2X1_322 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1261_), .B(_1227__bF_buf2), .Q(_1705_) );
NA3I1X1 NA3I1X1_39 ( .gnd!(gnd!), .vdd!(vdd!), .AN(_1223_), .B(_1695_), .C(_1705_), .Q(_1706_) );
NA2I1X1 NA2I1X1_46 ( .gnd!(gnd!), .vdd!(vdd!), .AN(_1293_), .B(_1227__bF_buf4), .Q(_1707_) );
ON211X1 ON211X1_50 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1230__bF_buf3), .B(_1250_), .C(_1239_), .D(_1226__bF_buf4), .Q(_1708_) );
ON21X1 ON21X1_221 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1269_), .B(_1226__bF_buf1), .C(_1223_), .Q(_1709_) );
AND2X2 AND2X2_13 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1709_), .B(_1221__bF_buf2), .Q(_1710_) );
AN32X1 AN32X1_2 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1222__bF_buf5), .B(_1707_), .C(_1708_), .D(_1710_), .E(_1706_), .Q(_1711_) );
NA2X1 NA2X1_323 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1288_), .B(_1307_), .Q(_1712_) );
MU2IX1 MU2IX1_62 ( .gnd!(gnd!), .vdd!(vdd!), .IN0(_1712_), .IN1(_1650_), .Q(_1713_), .S(_1240__bF_buf6) );
MU2IX1 MU2IX1_63 ( .gnd!(gnd!), .vdd!(vdd!), .IN0(_1548_), .IN1(_1713_), .Q(_1714_), .S(_1252__bF_buf4) );
MU2X1 MU2X1_189 ( .gnd!(gnd!), .vdd!(vdd!), .IN0(_1714_), .IN1(_1320_), .Q(_1715_), .S(_1226__bF_buf6) );
ON22X1 ON22X1_13 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1711_), .B(_866__bF_buf4), .C(_1400_), .D(_1715_), .Q(_1716_) );
ON21X1 ON21X1_222 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1048__bF_buf1), .B(_931__bF_buf4), .C(ALU_b_9_), .Q(_1717_) );
NA3I1X1 NA3I1X1_40 ( .gnd!(gnd!), .vdd!(vdd!), .AN(ALU_b_9_), .B(_1143__bF_buf3), .C(_1203__bF_buf1), .Q(_1718_) );
NA3I1X1 NA3I1X1_41 ( .gnd!(gnd!), .vdd!(vdd!), .AN(_1287_), .B(_1717_), .C(_1718_), .Q(_1719_) );
INX1 INX1_104 ( .gnd!(gnd!), .vdd!(vdd!), .A(ALU_b_9_), .Q(_1720_) );
ON21X1 ON21X1_223 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1048__bF_buf1), .B(_931__bF_buf4), .C(_1720_), .Q(_1721_) );
NA3I1X1 NA3I1X1_42 ( .gnd!(gnd!), .vdd!(vdd!), .AN(_1720_), .B(_1143__bF_buf3), .C(_1203__bF_buf1), .Q(_1722_) );
NA3I1X1 NA3I1X1_43 ( .gnd!(gnd!), .vdd!(vdd!), .AN(ALU_a_9_), .B(_1721_), .C(_1722_), .Q(_1723_) );
NA2X1 NA2X1_324 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1719_), .B(_1723_), .Q(_1724_) );
ON211X1 ON211X1_51 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1676_), .B(_1668_), .C(_1663_), .D(_1724_), .Q(_1725_) );
AN21X1 AN21X1_103 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1666_), .B(_1665_), .C(_1306_), .Q(_1726_) );
NO2X1 NO2X1_144 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1668_), .B(_1724_), .Q(_1727_) );
AN32X1 AN32X1_3 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1726_), .B(_1719_), .C(_1723_), .D(_1681_), .E(_1727_), .Q(_1728_) );
NA2X1 NA2X1_325 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1728_), .B(_1725_), .Q(_1729_) );
NA2X1 NA2X1_326 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1729_), .B(_952__bF_buf3), .Q(_1730_) );
ON211X1 ON211X1_52 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1716_), .B(_952__bF_buf1), .C(_909__bF_buf4), .D(_1730_), .Q(_1731_) );
AN22X1 AN22X1_29 ( .gnd!(gnd!), .vdd!(vdd!), .A(_866__bF_buf2), .B(_1524__bF_buf3), .C(_1731_), .D(_1704_), .Q(ALU_r_9_) );
NA2X1 NA2X1_327 ( .gnd!(gnd!), .vdd!(vdd!), .A(ALU_a_10_), .B(ALU_b_10_), .Q(_1732_) );
NO2X1 NO2X1_145 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1732_), .B(_1328__bF_buf4), .Q(_1733_) );
ON22X1 ON22X1_14 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1329__bF_buf2), .B(_888__bF_buf2), .C(ALU_a_10_), .D(ALU_b_10_), .Q(_1734_) );
ON22X1 ON22X1_15 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1733_), .B(_1734_), .C(_1526__bF_buf2), .D(_1732_), .Q(_1735_) );
NA2X1 NA2X1_328 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1735_), .B(_1525__bF_buf0), .Q(_1736_) );
NO2X1 NO2X1_146 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1252__bF_buf4), .B(_1586_), .Q(_1737_) );
AND2X2 AND2X2_14 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1393_), .B(_1375_), .Q(_1738_) );
MU2IX1 MU2IX1_64 ( .gnd!(gnd!), .vdd!(vdd!), .IN0(_1685_), .IN1(_1738_), .Q(_1739_), .S(_1233__bF_buf4) );
NO2X1 NO2X1_147 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1230__bF_buf1), .B(_1739_), .Q(_1740_) );
NO2X1 NO2X1_148 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1737_), .B(_1740_), .Q(_1741_) );
MU2IX1 MU2IX1_65 ( .gnd!(gnd!), .vdd!(vdd!), .IN0(_1741_), .IN1(_1404_), .Q(_1742_), .S(_1226__bF_buf5) );
NA2X1 NA2X1_329 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1362_), .B(_1227__bF_buf4), .Q(_1743_) );
AND2X2 AND2X2_15 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1743_), .B(_1223_), .Q(_1744_) );
NA2X1 NA2X1_330 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1365_), .B(_1227__bF_buf1), .Q(_1745_) );
AND3X4 AND3X4_3 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1745_), .B(ALU_func7_5_bF_buf0), .C(_1695_), .Q(_1746_) );
NO2X1 NO2X1_149 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1227__bF_buf6), .B(_1348_), .Q(_1747_) );
ON21X1 ON21X1_224 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1397_), .B(_1226__bF_buf3), .C(_1222__bF_buf4), .Q(_1748_) );
ON32X1 ON32X1_1 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1222__bF_buf4), .B(_1744_), .C(_1746_), .D(_1747_), .E(_1748_), .Q(_1749_) );
AO22X2 AO22X2_24 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1322__bF_buf2), .B(_1742_), .C(_1749_), .D(EXT_type_bF_buf2), .Q(_1750_) );
AN21X1 AN21X1_104 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1722_), .B(_1721_), .C(ALU_a_9_), .Q(_1751_) );
AN21X1 AN21X1_105 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1718_), .B(_1717_), .C(_1287_), .Q(_1752_) );
ON211X1 ON211X1_53 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1751_), .B(_1752_), .C(_1663_), .D(_1667_), .Q(_1753_) );
AN21X1 AN21X1_106 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1722_), .B(_1721_), .C(_1287_), .Q(_1754_) );
AN21X1 AN21X1_107 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1726_), .B(_1723_), .C(_1754_), .Q(_1755_) );
ON21X1 ON21X1_225 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1676_), .B(_1753_), .C(_1755_), .Q(_1756_) );
ON21X1 ON21X1_226 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1048__bF_buf3), .B(_931__bF_buf1), .C(ALU_b_10_), .Q(_1757_) );
NA3I1X1 NA3I1X1_44 ( .gnd!(gnd!), .vdd!(vdd!), .AN(ALU_b_10_), .B(_1143__bF_buf4), .C(_1203__bF_buf4), .Q(_1758_) );
NA3I1X1 NA3I1X1_45 ( .gnd!(gnd!), .vdd!(vdd!), .AN(ALU_a_10_), .B(_1757_), .C(_1758_), .Q(_1759_) );
INX1 INX1_105 ( .gnd!(gnd!), .vdd!(vdd!), .A(ALU_b_10_), .Q(_1760_) );
ON21X1 ON21X1_227 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1048__bF_buf0), .B(_931__bF_buf0), .C(_1760_), .Q(_1761_) );
NA3I1X1 NA3I1X1_46 ( .gnd!(gnd!), .vdd!(vdd!), .AN(_1760_), .B(_1143__bF_buf4), .C(_1203__bF_buf4), .Q(_1762_) );
NA3I1X1 NA3I1X1_47 ( .gnd!(gnd!), .vdd!(vdd!), .AN(_1289_), .B(_1761_), .C(_1762_), .Q(_1763_) );
NA2X1 NA2X1_331 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1763_), .B(_1759_), .Q(_1764_) );
NA2X1 NA2X1_332 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1756_), .B(_1764_), .Q(_1765_) );
NA2X1 NA2X1_333 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1681_), .B(_1727_), .Q(_1766_) );
NA3I1X1 NA3I1X1_48 ( .gnd!(gnd!), .vdd!(vdd!), .AN(_1764_), .B(_1755_), .C(_1766_), .Q(_1767_) );
NA2X1 NA2X1_334 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1765_), .B(_1767_), .Q(_1768_) );
NA2X1 NA2X1_335 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1768_), .B(_952__bF_buf4), .Q(_1769_) );
ON211X1 ON211X1_54 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1750_), .B(_952__bF_buf1), .C(_909__bF_buf4), .D(_1769_), .Q(_1770_) );
AN22X1 AN22X1_30 ( .gnd!(gnd!), .vdd!(vdd!), .A(_866__bF_buf5), .B(_1524__bF_buf1), .C(_1770_), .D(_1736_), .Q(ALU_r_10_) );
NA2X1 NA2X1_336 ( .gnd!(gnd!), .vdd!(vdd!), .A(ALU_a_11_), .B(ALU_b_11_), .Q(_1771_) );
NO2X1 NO2X1_150 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1771_), .B(_1328__bF_buf4), .Q(_1772_) );
ON22X1 ON22X1_16 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1329__bF_buf2), .B(_888__bF_buf2), .C(ALU_a_11_), .D(ALU_b_11_), .Q(_1773_) );
ON22X1 ON22X1_17 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1772_), .B(_1773_), .C(_1526__bF_buf2), .D(_1771_), .Q(_1774_) );
NA2X1 NA2X1_337 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1774_), .B(_1525__bF_buf3), .Q(_1775_) );
NA2X1 NA2X1_338 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1434_), .B(_1227__bF_buf4), .Q(_1776_) );
AND3X4 AND3X4_4 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1776_), .B(ALU_func7_5_bF_buf0), .C(_1695_), .Q(_1777_) );
NA2I1X1 NA2I1X1_47 ( .gnd!(gnd!), .vdd!(vdd!), .AN(_1438_), .B(_1227__bF_buf4), .Q(_1778_) );
AND2X2 AND2X2_16 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1778_), .B(_1223_), .Q(_1779_) );
NO2X1 NO2X1_151 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1226__bF_buf3), .B(_1444_), .Q(_1780_) );
ON211X1 ON211X1_55 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1230__bF_buf3), .B(_1429_), .C(_1428_), .D(_1226__bF_buf4), .Q(_1781_) );
NA2X1 NA2X1_339 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1781_), .B(_1222__bF_buf4), .Q(_1782_) );
ON32X1 ON32X1_2 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1222__bF_buf4), .B(_1777_), .C(_1779_), .D(_1780_), .E(_1782_), .Q(_1783_) );
NA2X1 NA2X1_340 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1283_), .B(_1290_), .Q(_1784_) );
MU2IX1 MU2IX1_66 ( .gnd!(gnd!), .vdd!(vdd!), .IN0(_1784_), .IN1(_1712_), .Q(_1785_), .S(_1240__bF_buf6) );
MU2IX1 MU2IX1_67 ( .gnd!(gnd!), .vdd!(vdd!), .IN0(_1651_), .IN1(_1785_), .Q(_1786_), .S(_1252__bF_buf4) );
MU2IX1 MU2IX1_68 ( .gnd!(gnd!), .vdd!(vdd!), .IN0(_1453_), .IN1(_1786_), .Q(_1787_), .S(_1227__bF_buf3) );
AO22X2 AO22X2_25 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1322__bF_buf0), .B(_1787_), .C(_1783_), .D(EXT_type_bF_buf6), .Q(_1788_) );
NA3I1X1 NA3I1X1_49 ( .gnd!(gnd!), .vdd!(vdd!), .AN(_1289_), .B(_1757_), .C(_1758_), .Q(_1789_) );
INX1 INX1_106 ( .gnd!(gnd!), .vdd!(vdd!), .A(ALU_b_11_), .Q(_1790_) );
ON21X1 ON21X1_228 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1048__bF_buf3), .B(_931__bF_buf1), .C(_1790_), .Q(_1791_) );
NA3I1X1 NA3I1X1_50 ( .gnd!(gnd!), .vdd!(vdd!), .AN(_1790_), .B(_1143__bF_buf2), .C(_1203__bF_buf4), .Q(_1792_) );
AN21X1 AN21X1_108 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1792_), .B(_1791_), .C(_1282_), .Q(_1793_) );
ON21X1 ON21X1_229 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1048__bF_buf3), .B(_931__bF_buf1), .C(ALU_b_11_), .Q(_1794_) );
NA3I1X1 NA3I1X1_51 ( .gnd!(gnd!), .vdd!(vdd!), .AN(ALU_b_11_), .B(_1143__bF_buf2), .C(_1203__bF_buf4), .Q(_1795_) );
AN21X1 AN21X1_109 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1795_), .B(_1794_), .C(ALU_a_11_), .Q(_1796_) );
NO2X1 NO2X1_152 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1793_), .B(_1796_), .Q(_1797_) );
NA3I1X1 NA3I1X1_52 ( .gnd!(gnd!), .vdd!(vdd!), .AN(_1797_), .B(_1789_), .C(_1765_), .Q(_1798_) );
NA2X1 NA2X1_341 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1765_), .B(_1789_), .Q(_1799_) );
NA2X1 NA2X1_342 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1799_), .B(_1797_), .Q(_1800_) );
NA2X1 NA2X1_343 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1800_), .B(_1798_), .Q(_1801_) );
NA2X1 NA2X1_344 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1801_), .B(_952__bF_buf2), .Q(_1802_) );
ON211X1 ON211X1_56 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1788_), .B(_952__bF_buf2), .C(_909__bF_buf4), .D(_1802_), .Q(_1803_) );
AN22X1 AN22X1_31 ( .gnd!(gnd!), .vdd!(vdd!), .A(_866__bF_buf3), .B(_1524__bF_buf2), .C(_1803_), .D(_1775_), .Q(ALU_r_11_) );
NA2X1 NA2X1_345 ( .gnd!(gnd!), .vdd!(vdd!), .A(ALU_a_12_), .B(ALU_b_12_), .Q(_1804_) );
NO2X1 NO2X1_153 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1804_), .B(_1328__bF_buf3), .Q(_1805_) );
ON22X1 ON22X1_18 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1329__bF_buf2), .B(_888__bF_buf2), .C(ALU_a_12_), .D(ALU_b_12_), .Q(_1806_) );
ON22X1 ON22X1_19 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1805_), .B(_1806_), .C(_1526__bF_buf0), .D(_1804_), .Q(_1807_) );
NA2X1 NA2X1_346 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1807_), .B(_1525__bF_buf1), .Q(_1808_) );
AN21X1 AN21X1_110 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1718_), .B(_1717_), .C(ALU_a_9_), .Q(_1809_) );
ON21X1 ON21X1_230 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1809_), .B(_1663_), .C(_1719_), .Q(_1810_) );
NA3I1X1 NA3I1X1_53 ( .gnd!(gnd!), .vdd!(vdd!), .AN(_1282_), .B(_1794_), .C(_1795_), .Q(_1811_) );
AN21X1 AN21X1_111 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1789_), .B(_1811_), .C(_1796_), .Q(_1812_) );
AN31X1 AN31X1_43 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1764_), .B(_1797_), .C(_1810_), .D(_1812_), .Q(_1813_) );
NA3I1X1 NA3I1X1_54 ( .gnd!(gnd!), .vdd!(vdd!), .AN(ALU_a_11_), .B(_1791_), .C(_1792_), .Q(_1814_) );
NA2X1 NA2X1_347 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1811_), .B(_1814_), .Q(_1815_) );
NA3I1X1 NA3I1X1_55 ( .gnd!(gnd!), .vdd!(vdd!), .AN(_1815_), .B(_1764_), .C(_1727_), .Q(_1816_) );
ON21X1 ON21X1_231 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1676_), .B(_1816_), .C(_1813_), .Q(_1817_) );
INX1 INX1_107 ( .gnd!(gnd!), .vdd!(vdd!), .A(ALU_b_12_), .Q(_1818_) );
ON21X1 ON21X1_232 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1048__bF_buf2), .B(_931__bF_buf0), .C(_1818_), .Q(_1819_) );
NA3I1X1 NA3I1X1_56 ( .gnd!(gnd!), .vdd!(vdd!), .AN(_1818_), .B(_1143__bF_buf4), .C(_1203__bF_buf2), .Q(_1820_) );
AN21X1 AN21X1_112 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1820_), .B(_1819_), .C(ALU_a_12_), .Q(_1821_) );
ON21X1 ON21X1_233 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1048__bF_buf0), .B(_931__bF_buf5), .C(ALU_b_12_), .Q(_1822_) );
NA3I1X1 NA3I1X1_57 ( .gnd!(gnd!), .vdd!(vdd!), .AN(ALU_b_12_), .B(_1143__bF_buf4), .C(_1203__bF_buf2), .Q(_1823_) );
AN21X1 AN21X1_113 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1823_), .B(_1822_), .C(_1284_), .Q(_1824_) );
NO2X1 NO2X1_154 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1821_), .B(_1824_), .Q(_1825_) );
NA2I1X1 NA2I1X1_48 ( .gnd!(gnd!), .vdd!(vdd!), .AN(_1825_), .B(_1817_), .Q(_1826_) );
ON211X1 ON211X1_57 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1676_), .B(_1816_), .C(_1813_), .D(_1825_), .Q(_1827_) );
NA2X1 NA2X1_348 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1826_), .B(_1827_), .Q(_1828_) );
NA2X1 NA2X1_349 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1828_), .B(_952__bF_buf3), .Q(_1829_) );
MU2IX1 MU2IX1_69 ( .gnd!(gnd!), .vdd!(vdd!), .IN0(_1507_), .IN1(_1498_), .Q(_1830_), .S(_1226__bF_buf0) );
NA2X1 NA2X1_350 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1830_), .B(_1222__bF_buf3), .Q(_1831_) );
NA2X1 NA2X1_351 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1500_), .B(_1227__bF_buf4), .Q(_1832_) );
AND2X2 AND2X2_17 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1433_), .B(_1695_), .Q(_1833_) );
ON211X1 ON211X1_58 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1223_), .B(_1833_), .C(_1832_), .D(_1221__bF_buf1), .Q(_1834_) );
AND2X2 AND2X2_18 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1517_), .B(_1226__bF_buf6), .Q(_1835_) );
NA2X1 NA2X1_352 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1686_), .B(_1230__bF_buf2), .Q(_1836_) );
AND2X2 AND2X2_19 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1390_), .B(_1394_), .Q(_1837_) );
MU2X1 MU2X1_190 ( .gnd!(gnd!), .vdd!(vdd!), .IN0(_1837_), .IN1(_1738_), .Q(_1838_), .S(_1240__bF_buf3) );
NA2X1 NA2X1_353 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1838_), .B(_1252__bF_buf2), .Q(_1839_) );
AN31X1 AN31X1_44 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1227__bF_buf5), .B(_1836_), .C(_1839_), .D(_1835_), .Q(_1840_) );
AO32X4 AO32X4_1 ( .gnd!(gnd!), .vdd!(vdd!), .A(EXT_type_bF_buf6), .B(_1831_), .C(_1834_), .D(_1840_), .E(_1322__bF_buf0), .Q(_1841_) );
ON211X1 ON211X1_59 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1841_), .B(_952__bF_buf1), .C(_909__bF_buf4), .D(_1829_), .Q(_1842_) );
AN22X1 AN22X1_32 ( .gnd!(gnd!), .vdd!(vdd!), .A(_866__bF_buf3), .B(_1524__bF_buf2), .C(_1842_), .D(_1808_), .Q(ALU_r_12_) );
NA2X1 NA2X1_354 ( .gnd!(gnd!), .vdd!(vdd!), .A(ALU_a_13_), .B(ALU_b_13_), .Q(_1843_) );
NO2X1 NO2X1_155 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1843_), .B(_1328__bF_buf3), .Q(_1844_) );
ON22X1 ON22X1_20 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1329__bF_buf2), .B(_888__bF_buf2), .C(ALU_a_13_), .D(ALU_b_13_), .Q(_1845_) );
ON22X1 ON22X1_21 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1844_), .B(_1845_), .C(_1526__bF_buf0), .D(_1843_), .Q(_1846_) );
NA2X1 NA2X1_355 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1846_), .B(_1525__bF_buf1), .Q(_1847_) );
NA3I1X1 NA3I1X1_58 ( .gnd!(gnd!), .vdd!(vdd!), .AN(_1284_), .B(_1822_), .C(_1823_), .Q(_1848_) );
ON21X1 ON21X1_234 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1048__bF_buf2), .B(_931__bF_buf0), .C(ALU_b_13_), .Q(_1849_) );
NA3I1X1 NA3I1X1_59 ( .gnd!(gnd!), .vdd!(vdd!), .AN(ALU_b_13_), .B(_1143__bF_buf4), .C(_1203__bF_buf2), .Q(_1850_) );
NA3I1X1 NA3I1X1_60 ( .gnd!(gnd!), .vdd!(vdd!), .AN(ALU_a_13_), .B(_1849_), .C(_1850_), .Q(_1851_) );
INX1 INX1_108 ( .gnd!(gnd!), .vdd!(vdd!), .A(ALU_b_13_), .Q(_1852_) );
ON21X1 ON21X1_235 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1048__bF_buf2), .B(_931__bF_buf0), .C(_1852_), .Q(_1853_) );
NA3I1X1 NA3I1X1_61 ( .gnd!(gnd!), .vdd!(vdd!), .AN(_1852_), .B(_1143__bF_buf4), .C(_1203__bF_buf2), .Q(_1854_) );
NA3I1X1 NA3I1X1_62 ( .gnd!(gnd!), .vdd!(vdd!), .AN(_1276_), .B(_1853_), .C(_1854_), .Q(_1855_) );
NA2X1 NA2X1_356 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1851_), .B(_1855_), .Q(_1856_) );
NA3I1X1 NA3I1X1_63 ( .gnd!(gnd!), .vdd!(vdd!), .AN(_1856_), .B(_1848_), .C(_1826_), .Q(_1857_) );
NA2X1 NA2X1_357 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1826_), .B(_1848_), .Q(_1858_) );
NA2X1 NA2X1_358 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1858_), .B(_1856_), .Q(_1859_) );
NA2X1 NA2X1_359 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1859_), .B(_1857_), .Q(_1860_) );
NA2X1 NA2X1_360 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1860_), .B(_952__bF_buf3), .Q(_1861_) );
ON21X1 ON21X1_236 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1538_), .B(_1226__bF_buf1), .C(_1833_), .Q(_1862_) );
NA2X1 NA2X1_361 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1535_), .B(_1227__bF_buf2), .Q(_1863_) );
NA2X1 NA2X1_362 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1863_), .B(_1223_), .Q(_1864_) );
ON211X1 ON211X1_60 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1862_), .B(_1223_), .C(_1864_), .D(_1221__bF_buf2), .Q(_1865_) );
AND3X4 AND3X4_5 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1532_), .B(_1533_), .C(_1226__bF_buf4), .Q(_1866_) );
AND2X2 AND2X2_20 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1544_), .B(_1227__bF_buf2), .Q(_1867_) );
ON31X1 ON31X1_40 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1221__bF_buf2), .B(_1866_), .C(_1867_), .D(_1865_), .Q(_1868_) );
NA2X1 NA2X1_363 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1277_), .B(_1285_), .Q(_1869_) );
MU2IX1 MU2IX1_70 ( .gnd!(gnd!), .vdd!(vdd!), .IN0(_1869_), .IN1(_1784_), .Q(_1870_), .S(_1240__bF_buf3) );
MU2X1 MU2X1_191 ( .gnd!(gnd!), .vdd!(vdd!), .IN0(_1870_), .IN1(_1713_), .Q(_1871_), .S(_1230__bF_buf2) );
NA2X1 NA2X1_364 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1871_), .B(_1227__bF_buf3), .Q(_1872_) );
ON21X1 ON21X1_237 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1227__bF_buf3), .B(_1549_), .C(_1872_), .Q(_1873_) );
AO22X2 AO22X2_26 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1322__bF_buf3), .B(_1873_), .C(_1868_), .D(EXT_type_bF_buf2), .Q(_1874_) );
ON211X1 ON211X1_61 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1874_), .B(_952__bF_buf2), .C(_1861_), .D(_909__bF_buf4), .Q(_1875_) );
AN22X1 AN22X1_33 ( .gnd!(gnd!), .vdd!(vdd!), .A(_866__bF_buf2), .B(_1524__bF_buf3), .C(_1875_), .D(_1847_), .Q(ALU_r_13_) );
NA2X1 NA2X1_365 ( .gnd!(gnd!), .vdd!(vdd!), .A(ALU_a_14_), .B(ALU_b_14_), .Q(_1876_) );
NO2X1 NO2X1_156 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1876_), .B(_1328__bF_buf4), .Q(_1877_) );
ON22X1 ON22X1_22 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1329__bF_buf2), .B(_888__bF_buf2), .C(ALU_a_14_), .D(ALU_b_14_), .Q(_1878_) );
ON22X1 ON22X1_23 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1877_), .B(_1878_), .C(_1526__bF_buf2), .D(_1876_), .Q(_1879_) );
NA2X1 NA2X1_366 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1879_), .B(_1525__bF_buf0), .Q(_1880_) );
ON21X1 ON21X1_238 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1048__bF_buf0), .B(_931__bF_buf5), .C(ALU_b_14_), .Q(_1881_) );
NA3I1X1 NA3I1X1_64 ( .gnd!(gnd!), .vdd!(vdd!), .AN(ALU_b_14_), .B(_1143__bF_buf0), .C(_1203__bF_buf3), .Q(_1882_) );
NA3I1X1 NA3I1X1_65 ( .gnd!(gnd!), .vdd!(vdd!), .AN(ALU_a_14_), .B(_1881_), .C(_1882_), .Q(_1883_) );
INX1 INX1_109 ( .gnd!(gnd!), .vdd!(vdd!), .A(ALU_b_14_), .Q(_1884_) );
ON21X1 ON21X1_239 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1048__bF_buf0), .B(_931__bF_buf5), .C(_1884_), .Q(_1885_) );
NA3I1X1 NA3I1X1_66 ( .gnd!(gnd!), .vdd!(vdd!), .AN(_1884_), .B(_1143__bF_buf0), .C(_1203__bF_buf3), .Q(_1886_) );
NA3I1X1 NA3I1X1_67 ( .gnd!(gnd!), .vdd!(vdd!), .AN(_1278_), .B(_1885_), .C(_1886_), .Q(_1887_) );
NA2X1 NA2X1_367 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1887_), .B(_1883_), .Q(_1888_) );
NA3I1X1 NA3I1X1_68 ( .gnd!(gnd!), .vdd!(vdd!), .AN(ALU_a_13_), .B(_1853_), .C(_1854_), .Q(_1889_) );
NA3I1X1 NA3I1X1_69 ( .gnd!(gnd!), .vdd!(vdd!), .AN(_1276_), .B(_1849_), .C(_1850_), .Q(_1890_) );
NA2X1 NA2X1_368 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1848_), .B(_1890_), .Q(_1891_) );
NA2X1 NA2X1_369 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1891_), .B(_1889_), .Q(_1892_) );
NA3I1X1 NA3I1X1_70 ( .gnd!(gnd!), .vdd!(vdd!), .AN(ALU_a_12_), .B(_1822_), .C(_1823_), .Q(_1893_) );
NA3I1X1 NA3I1X1_71 ( .gnd!(gnd!), .vdd!(vdd!), .AN(_1284_), .B(_1819_), .C(_1820_), .Q(_1894_) );
AN22X1 AN22X1_34 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1893_), .B(_1894_), .C(_1851_), .D(_1855_), .Q(_1895_) );
NA2X1 NA2X1_370 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1817_), .B(_1895_), .Q(_1896_) );
NA2X1 NA2X1_371 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1896_), .B(_1892_), .Q(_1897_) );
NA2X1 NA2X1_372 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1897_), .B(_1888_), .Q(_1898_) );
NA3I1X1 NA3I1X1_72 ( .gnd!(gnd!), .vdd!(vdd!), .AN(_1888_), .B(_1892_), .C(_1896_), .Q(_1899_) );
AND2X2 AND2X2_21 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1898_), .B(_1899_), .Q(_1900_) );
NA2I1X1 NA2I1X1_49 ( .gnd!(gnd!), .vdd!(vdd!), .AN(_1578_), .B(_1227__bF_buf1), .Q(_1901_) );
AN31X1 AN31X1_45 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1227__bF_buf1), .B(_1575_), .C(_1578_), .D(_1641_), .Q(_1902_) );
NO2X1 NO2X1_157 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1223_), .B(_1902_), .Q(_1903_) );
AN211X1 AN211X1_5 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1223_), .B(_1901_), .C(_1222__bF_buf1), .D(_1903_), .Q(_1904_) );
AND2X2 AND2X2_22 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1582_), .B(_1227__bF_buf6), .Q(_1905_) );
AN311X1 AN311X1_3 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1226__bF_buf2), .B(_1572_), .C(_1573_), .D(_1221__bF_buf4), .E(_1905_), .Q(_1906_) );
ON21X1 ON21X1_240 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1906_), .B(_1904_), .C(EXT_type_bF_buf1), .Q(_1907_) );
AND2X2 AND2X2_23 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1387_), .B(_1391_), .Q(_1908_) );
MU2IX1 MU2IX1_71 ( .gnd!(gnd!), .vdd!(vdd!), .IN0(_1837_), .IN1(_1908_), .Q(_1909_), .S(_1233__bF_buf4) );
MU2IX1 MU2IX1_72 ( .gnd!(gnd!), .vdd!(vdd!), .IN0(_1739_), .IN1(_1909_), .Q(_1910_), .S(_1252__bF_buf2) );
NA2X1 NA2X1_373 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1910_), .B(_1227__bF_buf5), .Q(_1911_) );
ON21X1 ON21X1_241 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1227__bF_buf5), .B(_1587_), .C(_1911_), .Q(_1912_) );
NA2X1 NA2X1_374 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1912_), .B(_1322__bF_buf1), .Q(_1913_) );
AN31X1 AN31X1_46 ( .gnd!(gnd!), .vdd!(vdd!), .A(_941__bF_buf3), .B(_1913_), .C(_1907_), .D(_1525__bF_buf2), .Q(_1914_) );
ON21X1 ON21X1_242 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1900_), .B(_941__bF_buf0), .C(_1914_), .Q(_1915_) );
AN22X1 AN22X1_35 ( .gnd!(gnd!), .vdd!(vdd!), .A(_866__bF_buf5), .B(_1524__bF_buf1), .C(_1915_), .D(_1880_), .Q(ALU_r_14_) );
NA2X1 NA2X1_375 ( .gnd!(gnd!), .vdd!(vdd!), .A(ALU_a_15_), .B(ALU_b_15_), .Q(_1916_) );
NO2X1 NO2X1_158 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1916_), .B(_1328__bF_buf1), .Q(_1917_) );
ON22X1 ON22X1_24 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1329__bF_buf0), .B(_888__bF_buf1), .C(ALU_a_15_), .D(ALU_b_15_), .Q(_1918_) );
ON22X1 ON22X1_25 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1917_), .B(_1918_), .C(_1526__bF_buf1), .D(_1916_), .Q(_1919_) );
NA2X1 NA2X1_376 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1919_), .B(_1525__bF_buf0), .Q(_1920_) );
AN21X1 AN21X1_114 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1886_), .B(_1885_), .C(_1278_), .Q(_1921_) );
INX1 INX1_110 ( .gnd!(gnd!), .vdd!(vdd!), .A(ALU_b_15_), .Q(_1922_) );
ON21X1 ON21X1_243 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1048__bF_buf0), .B(_931__bF_buf0), .C(_1922_), .Q(_1923_) );
NA3I1X1 NA3I1X1_73 ( .gnd!(gnd!), .vdd!(vdd!), .AN(_1922_), .B(_1143__bF_buf0), .C(_1203__bF_buf2), .Q(_1924_) );
AN21X1 AN21X1_115 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1924_), .B(_1923_), .C(_1273_), .Q(_1925_) );
ON21X1 ON21X1_244 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1048__bF_buf0), .B(_931__bF_buf0), .C(ALU_b_15_), .Q(_1926_) );
NA3I1X1 NA3I1X1_74 ( .gnd!(gnd!), .vdd!(vdd!), .AN(ALU_b_15_), .B(_1143__bF_buf0), .C(_1203__bF_buf2), .Q(_1927_) );
AN21X1 AN21X1_116 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1927_), .B(_1926_), .C(ALU_a_15_), .Q(_1928_) );
NO2X1 NO2X1_159 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1925_), .B(_1928_), .Q(_1929_) );
AN211X1 AN211X1_6 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1888_), .B(_1897_), .C(_1921_), .D(_1929_), .Q(_1930_) );
NA3I1X1 NA3I1X1_75 ( .gnd!(gnd!), .vdd!(vdd!), .AN(_1278_), .B(_1881_), .C(_1882_), .Q(_1931_) );
NA3I1X1 NA3I1X1_76 ( .gnd!(gnd!), .vdd!(vdd!), .AN(_1273_), .B(_1926_), .C(_1927_), .Q(_1932_) );
NA3I1X1 NA3I1X1_77 ( .gnd!(gnd!), .vdd!(vdd!), .AN(ALU_a_15_), .B(_1923_), .C(_1924_), .Q(_1933_) );
NA2X1 NA2X1_377 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1932_), .B(_1933_), .Q(_1934_) );
AN21X1 AN21X1_117 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1898_), .B(_1931_), .C(_1934_), .Q(_1935_) );
NO2X1 NO2X1_160 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1930_), .B(_1935_), .Q(_1936_) );
MU2IX1 MU2IX1_73 ( .gnd!(gnd!), .vdd!(vdd!), .IN0(_1646_), .IN1(_1635_), .Q(_1937_), .S(_1226__bF_buf4) );
NA2X1 NA2X1_378 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1937_), .B(_1222__bF_buf2), .Q(_1938_) );
NO2X1 NO2X1_161 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1223_), .B(_1265_), .Q(_1939_) );
INX1 INX1_111 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1939_), .Q(_1940_) );
NA2X1 NA2X1_379 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1221__bF_buf1), .B(_1940_), .Q(_1941_) );
NA2X1 NA2X1_380 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1941_), .B(EXT_type_bF_buf1), .Q(_1942_) );
NA2X1 NA2X1_381 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1637_), .B(_1227__bF_buf1), .Q(_1943_) );
ON31X1 ON31X1_41 ( .gnd!(gnd!), .vdd!(vdd!), .A(ALU_func7_5_bF_buf1), .B(_866__bF_buf1), .C(_1943_), .D(_1942_), .Q(_1944_) );
NA2X1 NA2X1_382 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1274_), .B(_1279_), .Q(_1945_) );
MU2IX1 MU2IX1_74 ( .gnd!(gnd!), .vdd!(vdd!), .IN0(_1945_), .IN1(_1869_), .Q(_1946_), .S(_1240__bF_buf3) );
MU2X1 MU2X1_192 ( .gnd!(gnd!), .vdd!(vdd!), .IN0(_1946_), .IN1(_1785_), .Q(_1947_), .S(_1230__bF_buf2) );
MU2X1 MU2X1_193 ( .gnd!(gnd!), .vdd!(vdd!), .IN0(_1652_), .IN1(_1947_), .Q(_1948_), .S(_1227__bF_buf5) );
AN22X1 AN22X1_36 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1322__bF_buf1), .B(_1948_), .C(_1938_), .D(_1944_), .Q(_1949_) );
NA2X1 NA2X1_383 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1949_), .B(_941__bF_buf3), .Q(_1950_) );
ON211X1 ON211X1_62 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1936_), .B(_941__bF_buf4), .C(_909__bF_buf1), .D(_1950_), .Q(_1951_) );
AN22X1 AN22X1_37 ( .gnd!(gnd!), .vdd!(vdd!), .A(_866__bF_buf5), .B(_1524__bF_buf1), .C(_1951_), .D(_1920_), .Q(ALU_r_15_) );
NA2X1 NA2X1_384 ( .gnd!(gnd!), .vdd!(vdd!), .A(ALU_a_16_), .B(ALU_b_16_), .Q(_1952_) );
NO2X1 NO2X1_162 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1952_), .B(_1328__bF_buf4), .Q(_1953_) );
ON22X1 ON22X1_26 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1329__bF_buf4), .B(_888__bF_buf2), .C(ALU_a_16_), .D(ALU_b_16_), .Q(_1954_) );
ON22X1 ON22X1_27 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1953_), .B(_1954_), .C(_1526__bF_buf0), .D(_1952_), .Q(_1955_) );
NA2X1 NA2X1_385 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1955_), .B(_1525__bF_buf3), .Q(_1956_) );
MU2IX1 MU2IX1_75 ( .gnd!(gnd!), .vdd!(vdd!), .IN0(_1693_), .IN1(_1690_), .Q(_1957_), .S(_1227__bF_buf6) );
AN21X1 AN21X1_118 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1957_), .B(_1222__bF_buf3), .C(_1942_), .Q(_1958_) );
NO2X1 NO2X1_163 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1226__bF_buf6), .B(_1684_), .Q(_1959_) );
NO2X1 NO2X1_164 ( .gnd!(gnd!), .vdd!(vdd!), .A(EXT_type_bF_buf6), .B(_1222__bF_buf2), .Q(_1960_) );
ON21X1 ON21X1_245 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1273_), .B(_1242__bF_buf0), .C(_1383_), .Q(_1961_) );
MU2IX1 MU2IX1_76 ( .gnd!(gnd!), .vdd!(vdd!), .IN0(_1908_), .IN1(_1961_), .Q(_1962_), .S(_1233__bF_buf4) );
NA2X1 NA2X1_386 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1962_), .B(_1252__bF_buf2), .Q(_1963_) );
ON21X1 ON21X1_246 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1838_), .B(_1252__bF_buf2), .C(_1963_), .Q(_1964_) );
NA2X1 NA2X1_387 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1964_), .B(_1227__bF_buf0), .Q(_1965_) );
NA2X1 NA2X1_388 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1687_), .B(_1226__bF_buf6), .Q(_1966_) );
AO32X4 AO32X4_2 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1322__bF_buf3), .B(_1965_), .C(_1966_), .D(_1959_), .E(_1960_), .Q(_1967_) );
AN21X1 AN21X1_119 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1762_), .B(_1761_), .C(ALU_a_10_), .Q(_1968_) );
AN21X1 AN21X1_120 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1758_), .B(_1757_), .C(_1289_), .Q(_1969_) );
ON211X1 ON211X1_63 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1968_), .B(_1969_), .C(_1811_), .D(_1814_), .Q(_1970_) );
ON211X1 ON211X1_64 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1821_), .B(_1824_), .C(_1890_), .D(_1889_), .Q(_1971_) );
AN21X1 AN21X1_121 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1886_), .B(_1885_), .C(ALU_a_14_), .Q(_1972_) );
AN21X1 AN21X1_122 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1882_), .B(_1881_), .C(_1278_), .Q(_1973_) );
ON211X1 ON211X1_65 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1972_), .B(_1973_), .C(_1932_), .D(_1933_), .Q(_1974_) );
NO2X1 NO2X1_165 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1971_), .B(_1974_), .Q(_1975_) );
NA3I1X1 NA3I1X1_78 ( .gnd!(gnd!), .vdd!(vdd!), .AN(_1970_), .B(_1727_), .C(_1975_), .Q(_1976_) );
AN21X1 AN21X1_123 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1762_), .B(_1761_), .C(_1289_), .Q(_1977_) );
NO2X1 NO2X1_166 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1977_), .B(_1793_), .Q(_1978_) );
ON22X1 ON22X1_28 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1970_), .B(_1755_), .C(_1978_), .D(_1796_), .Q(_1979_) );
NA2X1 NA2X1_389 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1921_), .B(_1933_), .Q(_1980_) );
ON211X1 ON211X1_66 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1892_), .B(_1974_), .C(_1932_), .D(_1980_), .Q(_1981_) );
AN21X1 AN21X1_124 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1979_), .B(_1975_), .C(_1981_), .Q(_1982_) );
ON21X1 ON21X1_247 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1676_), .B(_1976_), .C(_1982_), .Q(_1983_) );
INX1 INX1_112 ( .gnd!(gnd!), .vdd!(vdd!), .A(ALU_a_16_), .Q(_1984_) );
NA2X1 NA2X1_390 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1212__bF_buf4), .B(ALU_b_16_), .Q(_1985_) );
INX1 INX1_113 ( .gnd!(gnd!), .vdd!(vdd!), .A(ALU_b_16_), .Q(_1986_) );
NA2X1 NA2X1_391 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1059__bF_buf0), .B(_1986_), .Q(_1987_) );
NA3I1X1 NA3I1X1_79 ( .gnd!(gnd!), .vdd!(vdd!), .AN(_1984_), .B(_1985_), .C(_1987_), .Q(_1988_) );
NA2X1 NA2X1_392 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1212__bF_buf4), .B(_1986_), .Q(_1989_) );
NA2X1 NA2X1_393 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1059__bF_buf0), .B(ALU_b_16_), .Q(_1990_) );
NA3I1X1 NA3I1X1_80 ( .gnd!(gnd!), .vdd!(vdd!), .AN(ALU_a_16_), .B(_1989_), .C(_1990_), .Q(_1991_) );
AND2X2 AND2X2_24 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1988_), .B(_1991_), .Q(_1992_) );
NA2X1 NA2X1_394 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1983_), .B(_1992_), .Q(_1993_) );
NA3X1 NA3X1_4 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1888_), .B(_1929_), .C(_1895_), .Q(_1994_) );
NO2X1 NO2X1_167 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1994_), .B(_1816_), .Q(_1995_) );
AN21X1 AN21X1_125 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1850_), .B(_1849_), .C(ALU_a_13_), .Q(_1996_) );
ON21X1 ON21X1_248 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1996_), .B(_1848_), .C(_1890_), .Q(_1997_) );
ON21X1 ON21X1_249 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1928_), .B(_1931_), .C(_1932_), .Q(_1998_) );
AN31X1 AN31X1_47 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1888_), .B(_1929_), .C(_1997_), .D(_1998_), .Q(_1999_) );
ON21X1 ON21X1_250 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1813_), .B(_1994_), .C(_1999_), .Q(_2000_) );
AN21X1 AN21X1_126 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1681_), .B(_1995_), .C(_2000_), .Q(_2001_) );
NA2X1 NA2X1_395 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1988_), .B(_1991_), .Q(_2002_) );
NA2X1 NA2X1_396 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2001_), .B(_2002_), .Q(_2003_) );
NA2X1 NA2X1_397 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2003_), .B(_1993_), .Q(_2004_) );
NA2X1 NA2X1_398 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2004_), .B(_952__bF_buf3), .Q(_2005_) );
ON311X1 ON311X1_4 ( .gnd!(gnd!), .vdd!(vdd!), .A(_952__bF_buf5), .B(_1958_), .C(_1967_), .D(_909__bF_buf3), .E(_2005_), .Q(_2006_) );
AN22X1 AN22X1_38 ( .gnd!(gnd!), .vdd!(vdd!), .A(_866__bF_buf0), .B(_1524__bF_buf0), .C(_2006_), .D(_1956_), .Q(ALU_r_16_) );
AN21X1 AN21X1_127 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1990_), .B(_1989_), .C(_1984_), .Q(_2007_) );
INX1 INX1_114 ( .gnd!(gnd!), .vdd!(vdd!), .A(ALU_b_17_), .Q(_2008_) );
NA2X1 NA2X1_399 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1212__bF_buf4), .B(_2008_), .Q(_2009_) );
NA2X1 NA2X1_400 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1059__bF_buf0), .B(ALU_b_17_), .Q(_2010_) );
NA2X1 NA2X1_401 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2010_), .B(_2009_), .Q(_2011_) );
NA2X1 NA2X1_402 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2011_), .B(ALU_a_17_), .Q(_2012_) );
INX1 INX1_115 ( .gnd!(gnd!), .vdd!(vdd!), .A(ALU_a_17_), .Q(_2013_) );
NA2X1 NA2X1_403 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1212__bF_buf4), .B(ALU_b_17_), .Q(_2014_) );
NA2X1 NA2X1_404 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1059__bF_buf0), .B(_2008_), .Q(_2015_) );
NA2X1 NA2X1_405 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2015_), .B(_2014_), .Q(_2016_) );
NA2X1 NA2X1_406 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2016_), .B(_2013_), .Q(_2017_) );
NA2X1 NA2X1_407 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2012_), .B(_2017_), .Q(_2018_) );
NA3I1X1 NA3I1X1_81 ( .gnd!(gnd!), .vdd!(vdd!), .AN(_2007_), .B(_2018_), .C(_1993_), .Q(_2019_) );
NA2X1 NA2X1_408 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2011_), .B(_2013_), .Q(_2020_) );
NA2X1 NA2X1_409 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2016_), .B(ALU_a_17_), .Q(_2021_) );
NA2X1 NA2X1_410 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2020_), .B(_2021_), .Q(_2022_) );
NO2X1 NO2X1_168 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2002_), .B(_2018_), .Q(_2023_) );
AN22X1 AN22X1_39 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2007_), .B(_2022_), .C(_1983_), .D(_2023_), .Q(_2024_) );
NA3I1X1 NA3I1X1_82 ( .gnd!(gnd!), .vdd!(vdd!), .AN(_941__bF_buf1), .B(_2024_), .C(_2019_), .Q(_2025_) );
MU2IX1 MU2IX1_77 ( .gnd!(gnd!), .vdd!(vdd!), .IN0(ALU_a_17_), .IN1(ALU_a_16_), .Q(_2026_), .S(_1235__bF_buf2) );
MU2IX1 MU2IX1_78 ( .gnd!(gnd!), .vdd!(vdd!), .IN0(_2026_), .IN1(_1945_), .Q(_2027_), .S(_1240__bF_buf3) );
MU2IX1 MU2IX1_79 ( .gnd!(gnd!), .vdd!(vdd!), .IN0(_2027_), .IN1(_1870_), .Q(_2028_), .S(_1230__bF_buf1) );
MU2IX1 MU2IX1_80 ( .gnd!(gnd!), .vdd!(vdd!), .IN0(_1714_), .IN1(_2028_), .Q(_2029_), .S(_1227__bF_buf3) );
MU2IX1 MU2IX1_81 ( .gnd!(gnd!), .vdd!(vdd!), .IN0(_2029_), .IN1(_1321_), .Q(_2030_), .S(_1221__bF_buf3) );
NA2X1 NA2X1_411 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2030_), .B(_866__bF_buf4), .Q(_2031_) );
NA2X1 NA2X1_412 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1262_), .B(_1222__bF_buf5), .Q(_2032_) );
NA2X1 NA2X1_413 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1941_), .B(ALU_func7_5_bF_buf2), .Q(_2033_) );
INX1 INX1_116 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2033_), .Q(_2034_) );
NA2X1 NA2X1_414 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2032_), .B(_2034_), .Q(_2035_) );
NA2X1 NA2X1_415 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1222__bF_buf1), .B(_1223_), .Q(_2036_) );
ON211X1 ON211X1_67 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1271_), .B(_2036_), .C(_2035_), .D(EXT_type_bF_buf4), .Q(_689_) );
AN31X1 AN31X1_48 ( .gnd!(gnd!), .vdd!(vdd!), .A(_941__bF_buf3), .B(_2031_), .C(_689_), .D(_1525__bF_buf2), .Q(_690_) );
ON22X1 ON22X1_29 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1329__bF_buf0), .B(_888__bF_buf3), .C(ALU_a_17_), .D(ALU_b_17_), .Q(_691_) );
AN31X1 AN31X1_49 ( .gnd!(gnd!), .vdd!(vdd!), .A(ALU_a_17_), .B(ALU_b_17_), .C(_1327_), .D(_691_), .Q(_692_) );
AN31X1 AN31X1_50 ( .gnd!(gnd!), .vdd!(vdd!), .A(ALU_a_17_), .B(ALU_b_17_), .C(_1330_), .D(_692_), .Q(_693_) );
AN221X1 AN221X1_5 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1525__bF_buf0), .B(_693_), .C(_690_), .D(_2025_), .E(_931__bF_buf3), .Q(ALU_r_17_) );
NA2X1 NA2X1_416 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1992_), .B(_2022_), .Q(_694_) );
NO2X1 NO2X1_169 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2013_), .B(_2016_), .Q(_695_) );
AN21X1 AN21X1_128 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2007_), .B(_2017_), .C(_695_), .Q(_696_) );
ON21X1 ON21X1_251 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2001_), .B(_694_), .C(_696_), .Q(_697_) );
INX1 INX1_117 ( .gnd!(gnd!), .vdd!(vdd!), .A(ALU_a_18_), .Q(_698_) );
EN3X1 EN3X1_3 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1212__bF_buf0), .B(_698_), .C(ALU_b_18_), .Q(_699_) );
NA2X1 NA2X1_417 ( .gnd!(gnd!), .vdd!(vdd!), .A(_697_), .B(_699_), .Q(_700_) );
EN3X1 EN3X1_4 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1212__bF_buf0), .B(ALU_a_18_), .C(ALU_b_18_), .Q(_701_) );
NA3I1X1 NA3I1X1_83 ( .gnd!(gnd!), .vdd!(vdd!), .AN(_695_), .B(_701_), .C(_2024_), .Q(_702_) );
NA3I1X1 NA3I1X1_84 ( .gnd!(gnd!), .vdd!(vdd!), .AN(_941__bF_buf1), .B(_700_), .C(_702_), .Q(_703_) );
NA2X1 NA2X1_418 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1344_), .B(_1384_), .Q(_704_) );
MU2IX1 MU2IX1_82 ( .gnd!(gnd!), .vdd!(vdd!), .IN0(_704_), .IN1(_1961_), .Q(_705_), .S(_1240__bF_buf4) );
MU2X1 MU2X1_194 ( .gnd!(gnd!), .vdd!(vdd!), .IN0(_1909_), .IN1(_705_), .Q(_706_), .S(_1252__bF_buf2) );
AND2X2 AND2X2_25 ( .gnd!(gnd!), .vdd!(vdd!), .A(_706_), .B(_1227__bF_buf3), .Q(_707_) );
ON31X1 ON31X1_42 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1227__bF_buf5), .B(_1737_), .C(_1740_), .D(_1222__bF_buf2), .Q(_708_) );
ON32X1 ON32X1_3 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1222__bF_buf2), .B(_1226__bF_buf5), .C(_1404_), .D(_708_), .E(_707_), .Q(_709_) );
NA2X1 NA2X1_419 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1366_), .B(_1222__bF_buf1), .Q(_710_) );
NA2X1 NA2X1_420 ( .gnd!(gnd!), .vdd!(vdd!), .A(_710_), .B(_2034_), .Q(_711_) );
INX1 INX1_118 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2036_), .Q(_712_) );
NA2X1 NA2X1_421 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1363_), .B(_712_), .Q(_713_) );
AN31X1 AN31X1_51 ( .gnd!(gnd!), .vdd!(vdd!), .A(EXT_type_bF_buf1), .B(_713_), .C(_711_), .D(_952__bF_buf0), .Q(_714_) );
ON21X1 ON21X1_252 ( .gnd!(gnd!), .vdd!(vdd!), .A(EXT_type_bF_buf2), .B(_709_), .C(_714_), .Q(_715_) );
INX1 INX1_119 ( .gnd!(gnd!), .vdd!(vdd!), .A(ALU_b_18_), .Q(_716_) );
AN21X1 AN21X1_129 ( .gnd!(gnd!), .vdd!(vdd!), .A(_698_), .B(_716_), .C(_1330_), .Q(_717_) );
ON31X1 ON31X1_43 ( .gnd!(gnd!), .vdd!(vdd!), .A(_698_), .B(_716_), .C(_1328__bF_buf0), .D(_717_), .Q(_718_) );
ON31X1 ON31X1_44 ( .gnd!(gnd!), .vdd!(vdd!), .A(_698_), .B(_716_), .C(_1526__bF_buf3), .D(_718_), .Q(_719_) );
ON21X1 ON21X1_253 ( .gnd!(gnd!), .vdd!(vdd!), .A(_719_), .B(_909__bF_buf2), .C(_1143__bF_buf1), .Q(_720_) );
AN31X1 AN31X1_52 ( .gnd!(gnd!), .vdd!(vdd!), .A(_909__bF_buf2), .B(_703_), .C(_715_), .D(_720_), .Q(ALU_r_18_) );
NA2X1 NA2X1_422 ( .gnd!(gnd!), .vdd!(vdd!), .A(ALU_a_19_), .B(ALU_b_19_), .Q(_721_) );
NO2X1 NO2X1_170 ( .gnd!(gnd!), .vdd!(vdd!), .A(_721_), .B(_1328__bF_buf1), .Q(_722_) );
ON22X1 ON22X1_30 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1329__bF_buf3), .B(_888__bF_buf3), .C(ALU_a_19_), .D(ALU_b_19_), .Q(_723_) );
ON22X1 ON22X1_31 ( .gnd!(gnd!), .vdd!(vdd!), .A(_722_), .B(_723_), .C(_1526__bF_buf1), .D(_721_), .Q(_724_) );
NA2X1 NA2X1_423 ( .gnd!(gnd!), .vdd!(vdd!), .A(_724_), .B(_1525__bF_buf3), .Q(_725_) );
NA2X1 NA2X1_424 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1212__bF_buf0), .B(_716_), .Q(_726_) );
NA2X1 NA2X1_425 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1059__bF_buf1), .B(ALU_b_18_), .Q(_727_) );
NA2X1 NA2X1_426 ( .gnd!(gnd!), .vdd!(vdd!), .A(_727_), .B(_726_), .Q(_728_) );
NA2X1 NA2X1_427 ( .gnd!(gnd!), .vdd!(vdd!), .A(_728_), .B(ALU_a_18_), .Q(_729_) );
INX1 INX1_120 ( .gnd!(gnd!), .vdd!(vdd!), .A(_729_), .Q(_730_) );
NA2X1 NA2X1_428 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1212__bF_buf1), .B(ALU_b_19_), .Q(_731_) );
INX1 INX1_121 ( .gnd!(gnd!), .vdd!(vdd!), .A(ALU_b_19_), .Q(_732_) );
NA2X1 NA2X1_429 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1059__bF_buf3), .B(_732_), .Q(_733_) );
NA3X1 NA3X1_5 ( .gnd!(gnd!), .vdd!(vdd!), .A(ALU_a_19_), .B(_731_), .C(_733_), .Q(_734_) );
NA2X1 NA2X1_430 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1212__bF_buf4), .B(_732_), .Q(_735_) );
NA2X1 NA2X1_431 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1059__bF_buf1), .B(ALU_b_19_), .Q(_736_) );
NA3I1X1 NA3I1X1_85 ( .gnd!(gnd!), .vdd!(vdd!), .AN(ALU_a_19_), .B(_735_), .C(_736_), .Q(_737_) );
AND2X2 AND2X2_26 ( .gnd!(gnd!), .vdd!(vdd!), .A(_734_), .B(_737_), .Q(_738_) );
AN211X1 AN211X1_7 ( .gnd!(gnd!), .vdd!(vdd!), .A(_699_), .B(_697_), .C(_730_), .D(_738_), .Q(_739_) );
NA2X1 NA2X1_432 ( .gnd!(gnd!), .vdd!(vdd!), .A(_734_), .B(_737_), .Q(_740_) );
AN21X1 AN21X1_130 ( .gnd!(gnd!), .vdd!(vdd!), .A(_700_), .B(_729_), .C(_740_), .Q(_741_) );
NO2X1 NO2X1_171 ( .gnd!(gnd!), .vdd!(vdd!), .A(_739_), .B(_741_), .Q(_742_) );
AND2X2 AND2X2_27 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1243_), .B(_1247_), .Q(_743_) );
MU2IX1 MU2IX1_83 ( .gnd!(gnd!), .vdd!(vdd!), .IN0(_743_), .IN1(_2026_), .Q(_744_), .S(_1240__bF_buf4) );
MU2IX1 MU2IX1_84 ( .gnd!(gnd!), .vdd!(vdd!), .IN0(_744_), .IN1(_1946_), .Q(_745_), .S(_1230__bF_buf1) );
MU2X1 MU2X1_195 ( .gnd!(gnd!), .vdd!(vdd!), .IN0(_745_), .IN1(_1786_), .Q(_746_), .S(_1226__bF_buf6) );
MU2IX1 MU2IX1_85 ( .gnd!(gnd!), .vdd!(vdd!), .IN0(_746_), .IN1(_1454_), .Q(_747_), .S(_1221__bF_buf3) );
AND2X2 AND2X2_28 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1435_), .B(_1222__bF_buf1), .Q(_748_) );
ON22X1 ON22X1_32 ( .gnd!(gnd!), .vdd!(vdd!), .A(_748_), .B(_2033_), .C(_1440_), .D(_2036_), .Q(_749_) );
MU2IX1 MU2IX1_86 ( .gnd!(gnd!), .vdd!(vdd!), .IN0(_749_), .IN1(_747_), .Q(_750_), .S(_866__bF_buf4) );
NA2X1 NA2X1_433 ( .gnd!(gnd!), .vdd!(vdd!), .A(_750_), .B(_941__bF_buf4), .Q(_751_) );
ON211X1 ON211X1_68 ( .gnd!(gnd!), .vdd!(vdd!), .A(_941__bF_buf4), .B(_742_), .C(_751_), .D(_909__bF_buf3), .Q(_752_) );
AN22X1 AN22X1_40 ( .gnd!(gnd!), .vdd!(vdd!), .A(_866__bF_buf3), .B(_1524__bF_buf2), .C(_752_), .D(_725_), .Q(ALU_r_19_) );
NA2X1 NA2X1_434 ( .gnd!(gnd!), .vdd!(vdd!), .A(ALU_a_20_), .B(ALU_b_20_), .Q(_753_) );
NO2X1 NO2X1_172 ( .gnd!(gnd!), .vdd!(vdd!), .A(_753_), .B(_1328__bF_buf1), .Q(_754_) );
ON22X1 ON22X1_33 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1329__bF_buf3), .B(_888__bF_buf3), .C(ALU_a_20_), .D(ALU_b_20_), .Q(_755_) );
ON22X1 ON22X1_34 ( .gnd!(gnd!), .vdd!(vdd!), .A(_754_), .B(_755_), .C(_1526__bF_buf1), .D(_753_), .Q(_756_) );
NA2X1 NA2X1_435 ( .gnd!(gnd!), .vdd!(vdd!), .A(_756_), .B(_1525__bF_buf1), .Q(_757_) );
NO2X1 NO2X1_173 ( .gnd!(gnd!), .vdd!(vdd!), .A(ALU_a_17_), .B(_2011_), .Q(_758_) );
ON21X1 ON21X1_254 ( .gnd!(gnd!), .vdd!(vdd!), .A(_758_), .B(_1988_), .C(_2012_), .Q(_759_) );
NA2X1 NA2X1_436 ( .gnd!(gnd!), .vdd!(vdd!), .A(_729_), .B(_734_), .Q(_760_) );
NO2X1 NO2X1_174 ( .gnd!(gnd!), .vdd!(vdd!), .A(_701_), .B(_740_), .Q(_761_) );
AN22X1 AN22X1_41 ( .gnd!(gnd!), .vdd!(vdd!), .A(_737_), .B(_760_), .C(_759_), .D(_761_), .Q(_762_) );
NA2X1 NA2X1_437 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2023_), .B(_761_), .Q(_763_) );
ON21X1 ON21X1_255 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2001_), .B(_763_), .C(_762_), .Q(_764_) );
INX1 INX1_122 ( .gnd!(gnd!), .vdd!(vdd!), .A(ALU_a_20_), .Q(_765_) );
NA2X1 NA2X1_438 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1212__bF_buf2), .B(ALU_b_20_), .Q(_766_) );
NA2I1X1 NA2I1X1_50 ( .gnd!(gnd!), .vdd!(vdd!), .AN(ALU_b_20_), .B(_1059__bF_buf1), .Q(_767_) );
NA3I1X1 NA3I1X1_86 ( .gnd!(gnd!), .vdd!(vdd!), .AN(_765_), .B(_766_), .C(_767_), .Q(_768_) );
NA2X1 NA2X1_439 ( .gnd!(gnd!), .vdd!(vdd!), .A(_767_), .B(_766_), .Q(_769_) );
NA2X1 NA2X1_440 ( .gnd!(gnd!), .vdd!(vdd!), .A(_769_), .B(_765_), .Q(_770_) );
NA2X1 NA2X1_441 ( .gnd!(gnd!), .vdd!(vdd!), .A(_770_), .B(_768_), .Q(_771_) );
NA2I1X1 NA2I1X1_51 ( .gnd!(gnd!), .vdd!(vdd!), .AN(_771_), .B(_764_), .Q(_772_) );
NA2I1X1 NA2I1X1_52 ( .gnd!(gnd!), .vdd!(vdd!), .AN(_764_), .B(_771_), .Q(_773_) );
AND2X2 AND2X2_29 ( .gnd!(gnd!), .vdd!(vdd!), .A(_773_), .B(_772_), .Q(_774_) );
NA2X1 NA2X1_442 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1341_), .B(_1345_), .Q(_775_) );
MU2IX1 MU2IX1_87 ( .gnd!(gnd!), .vdd!(vdd!), .IN0(_775_), .IN1(_704_), .Q(_776_), .S(_1240__bF_buf4) );
MU2X1 MU2X1_196 ( .gnd!(gnd!), .vdd!(vdd!), .IN0(_1962_), .IN1(_776_), .Q(_777_), .S(_1252__bF_buf2) );
NA2X1 NA2X1_443 ( .gnd!(gnd!), .vdd!(vdd!), .A(_777_), .B(_1227__bF_buf3), .Q(_778_) );
AN31X1 AN31X1_53 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1226__bF_buf6), .B(_1836_), .C(_1839_), .D(_1221__bF_buf0), .Q(_779_) );
AN22X1 AN22X1_42 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1518_), .B(_1221__bF_buf0), .C(_778_), .D(_779_), .Q(_780_) );
NA2I1X1 NA2I1X1_53 ( .gnd!(gnd!), .vdd!(vdd!), .AN(_780_), .B(_866__bF_buf4), .Q(_781_) );
AND2X2 AND2X2_30 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1501_), .B(_1222__bF_buf4), .Q(_782_) );
ON22X1 ON22X1_35 ( .gnd!(gnd!), .vdd!(vdd!), .A(_782_), .B(_2033_), .C(_1502_), .D(_2036_), .Q(_783_) );
NA2X1 NA2X1_444 ( .gnd!(gnd!), .vdd!(vdd!), .A(_783_), .B(EXT_type_bF_buf6), .Q(_784_) );
AN31X1 AN31X1_54 ( .gnd!(gnd!), .vdd!(vdd!), .A(_941__bF_buf3), .B(_781_), .C(_784_), .D(_1525__bF_buf2), .Q(_785_) );
ON21X1 ON21X1_256 ( .gnd!(gnd!), .vdd!(vdd!), .A(_941__bF_buf0), .B(_774_), .C(_785_), .Q(_786_) );
AN22X1 AN22X1_43 ( .gnd!(gnd!), .vdd!(vdd!), .A(_866__bF_buf2), .B(_1524__bF_buf3), .C(_786_), .D(_757_), .Q(ALU_r_20_) );
NA2X1 NA2X1_445 ( .gnd!(gnd!), .vdd!(vdd!), .A(ALU_a_21_), .B(ALU_b_21_), .Q(_787_) );
NO2X1 NO2X1_175 ( .gnd!(gnd!), .vdd!(vdd!), .A(_787_), .B(_1328__bF_buf1), .Q(_788_) );
ON22X1 ON22X1_36 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1329__bF_buf3), .B(_888__bF_buf1), .C(ALU_a_21_), .D(ALU_b_21_), .Q(_789_) );
ON22X1 ON22X1_37 ( .gnd!(gnd!), .vdd!(vdd!), .A(_788_), .B(_789_), .C(_1526__bF_buf1), .D(_787_), .Q(_790_) );
NA2X1 NA2X1_446 ( .gnd!(gnd!), .vdd!(vdd!), .A(_790_), .B(_1525__bF_buf4), .Q(_791_) );
INX1 INX1_123 ( .gnd!(gnd!), .vdd!(vdd!), .A(_768_), .Q(_792_) );
NO2I1X1 NO2I1X1_35 ( .gnd!(gnd!), .vdd!(vdd!), .AN(_761_), .B(_694_), .Q(_793_) );
NA2X1 NA2X1_447 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1983_), .B(_793_), .Q(_794_) );
NA3I1X1 NA3I1X1_87 ( .gnd!(gnd!), .vdd!(vdd!), .AN(ALU_a_20_), .B(_766_), .C(_767_), .Q(_795_) );
NA2X1 NA2X1_448 ( .gnd!(gnd!), .vdd!(vdd!), .A(_769_), .B(ALU_a_20_), .Q(_796_) );
AN22X1 AN22X1_44 ( .gnd!(gnd!), .vdd!(vdd!), .A(_795_), .B(_796_), .C(_794_), .D(_762_), .Q(_797_) );
NA2X1 NA2X1_449 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1212__bF_buf2), .B(ALU_b_21_), .Q(_798_) );
INX1 INX1_124 ( .gnd!(gnd!), .vdd!(vdd!), .A(ALU_b_21_), .Q(_799_) );
NA2X1 NA2X1_450 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1059__bF_buf1), .B(_799_), .Q(_800_) );
NA3X1 NA3X1_6 ( .gnd!(gnd!), .vdd!(vdd!), .A(ALU_a_21_), .B(_798_), .C(_800_), .Q(_801_) );
NA2X1 NA2X1_451 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1212__bF_buf2), .B(_799_), .Q(_802_) );
NA2X1 NA2X1_452 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1059__bF_buf2), .B(ALU_b_21_), .Q(_803_) );
NA3I1X1 NA3I1X1_88 ( .gnd!(gnd!), .vdd!(vdd!), .AN(ALU_a_21_), .B(_802_), .C(_803_), .Q(_804_) );
NA2X1 NA2X1_453 ( .gnd!(gnd!), .vdd!(vdd!), .A(_801_), .B(_804_), .Q(_805_) );
ON21X1 ON21X1_257 ( .gnd!(gnd!), .vdd!(vdd!), .A(_797_), .B(_792_), .C(_805_), .Q(_806_) );
NA3I1X1 NA3I1X1_89 ( .gnd!(gnd!), .vdd!(vdd!), .AN(_805_), .B(_768_), .C(_772_), .Q(_807_) );
NA2X1 NA2X1_454 ( .gnd!(gnd!), .vdd!(vdd!), .A(_806_), .B(_807_), .Q(_808_) );
NA2I1X1 NA2I1X1_54 ( .gnd!(gnd!), .vdd!(vdd!), .AN(_1871_), .B(_1226__bF_buf5), .Q(_809_) );
MU2IX1 MU2IX1_88 ( .gnd!(gnd!), .vdd!(vdd!), .IN0(ALU_a_21_), .IN1(ALU_a_20_), .Q(_810_), .S(_1235__bF_buf3) );
MU2IX1 MU2IX1_89 ( .gnd!(gnd!), .vdd!(vdd!), .IN0(_743_), .IN1(_810_), .Q(_811_), .S(_1233__bF_buf3) );
MU2IX1 MU2IX1_90 ( .gnd!(gnd!), .vdd!(vdd!), .IN0(_811_), .IN1(_2027_), .Q(_812_), .S(_1230__bF_buf1) );
AN21X1 AN21X1_131 ( .gnd!(gnd!), .vdd!(vdd!), .A(_812_), .B(_1227__bF_buf5), .C(_1221__bF_buf3), .Q(_813_) );
AO22X2 AO22X2_27 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1550_), .B(_1221__bF_buf3), .C(_809_), .D(_813_), .Q(_814_) );
NO2X1 NO2X1_176 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1221__bF_buf2), .B(_1539_), .Q(_815_) );
ON32X1 ON32X1_4 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1534_), .B(_1536_), .C(_2036_), .D(_2033_), .E(_815_), .Q(_816_) );
MU2IX1 MU2IX1_91 ( .gnd!(gnd!), .vdd!(vdd!), .IN0(_816_), .IN1(_814_), .Q(_817_), .S(_866__bF_buf4) );
NA2X1 NA2X1_455 ( .gnd!(gnd!), .vdd!(vdd!), .A(_817_), .B(_941__bF_buf2), .Q(_818_) );
ON211X1 ON211X1_69 ( .gnd!(gnd!), .vdd!(vdd!), .A(_941__bF_buf2), .B(_808_), .C(_818_), .D(_909__bF_buf3), .Q(_819_) );
AN22X1 AN22X1_45 ( .gnd!(gnd!), .vdd!(vdd!), .A(_866__bF_buf0), .B(_1524__bF_buf0), .C(_819_), .D(_791_), .Q(ALU_r_21_) );
NA2X1 NA2X1_456 ( .gnd!(gnd!), .vdd!(vdd!), .A(ALU_a_22_), .B(ALU_b_22_), .Q(_820_) );
NO2X1 NO2X1_177 ( .gnd!(gnd!), .vdd!(vdd!), .A(_820_), .B(_1328__bF_buf1), .Q(_821_) );
ON22X1 ON22X1_38 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1329__bF_buf0), .B(_888__bF_buf3), .C(ALU_a_22_), .D(ALU_b_22_), .Q(_822_) );
ON22X1 ON22X1_39 ( .gnd!(gnd!), .vdd!(vdd!), .A(_821_), .B(_822_), .C(_1526__bF_buf4), .D(_820_), .Q(_823_) );
NA2X1 NA2X1_457 ( .gnd!(gnd!), .vdd!(vdd!), .A(_823_), .B(_1525__bF_buf4), .Q(_824_) );
AN21X1 AN21X1_132 ( .gnd!(gnd!), .vdd!(vdd!), .A(_795_), .B(_796_), .C(_805_), .Q(_825_) );
NA2X1 NA2X1_458 ( .gnd!(gnd!), .vdd!(vdd!), .A(_764_), .B(_825_), .Q(_826_) );
NA2X1 NA2X1_459 ( .gnd!(gnd!), .vdd!(vdd!), .A(_768_), .B(_801_), .Q(_827_) );
NA2X1 NA2X1_460 ( .gnd!(gnd!), .vdd!(vdd!), .A(_827_), .B(_804_), .Q(_828_) );
INX1 INX1_125 ( .gnd!(gnd!), .vdd!(vdd!), .A(ALU_b_22_), .Q(_829_) );
NA2X1 NA2X1_461 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1212__bF_buf1), .B(_829_), .Q(_830_) );
NA2X1 NA2X1_462 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1059__bF_buf3), .B(ALU_b_22_), .Q(_831_) );
AN21X1 AN21X1_133 ( .gnd!(gnd!), .vdd!(vdd!), .A(_831_), .B(_830_), .C(ALU_a_22_), .Q(_832_) );
INX1 INX1_126 ( .gnd!(gnd!), .vdd!(vdd!), .A(_832_), .Q(_833_) );
INX1 INX1_127 ( .gnd!(gnd!), .vdd!(vdd!), .A(ALU_a_22_), .Q(_835_) );
NA2X1 NA2X1_463 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1212__bF_buf1), .B(ALU_b_22_), .Q(_836_) );
NA2X1 NA2X1_464 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1059__bF_buf3), .B(_829_), .Q(_837_) );
AN21X1 AN21X1_134 ( .gnd!(gnd!), .vdd!(vdd!), .A(_837_), .B(_836_), .C(_835_), .Q(_838_) );
INX1 INX1_128 ( .gnd!(gnd!), .vdd!(vdd!), .A(_838_), .Q(_839_) );
AN22X1 AN22X1_46 ( .gnd!(gnd!), .vdd!(vdd!), .A(_833_), .B(_839_), .C(_826_), .D(_828_), .Q(_840_) );
NA2X1 NA2X1_465 ( .gnd!(gnd!), .vdd!(vdd!), .A(_839_), .B(_833_), .Q(_841_) );
AN221X1 AN221X1_6 ( .gnd!(gnd!), .vdd!(vdd!), .A(_804_), .B(_827_), .C(_764_), .D(_825_), .E(_841_), .Q(_842_) );
ON21X1 ON21X1_258 ( .gnd!(gnd!), .vdd!(vdd!), .A(_840_), .B(_842_), .C(_952__bF_buf3), .Q(_843_) );
NO2X1 NO2X1_178 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1226__bF_buf2), .B(_1587_), .Q(_844_) );
NA2X1 NA2X1_466 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1337_), .B(_1342_), .Q(_845_) );
MU2X1 MU2X1_197 ( .gnd!(gnd!), .vdd!(vdd!), .IN0(_845_), .IN1(_775_), .Q(_846_), .S(_1240__bF_buf2) );
NA2X1 NA2X1_467 ( .gnd!(gnd!), .vdd!(vdd!), .A(_846_), .B(_1252__bF_buf0), .Q(_847_) );
ON21X1 ON21X1_259 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1252__bF_buf2), .B(_705_), .C(_847_), .Q(_848_) );
MU2X1 MU2X1_198 ( .gnd!(gnd!), .vdd!(vdd!), .IN0(_848_), .IN1(_1910_), .Q(_849_), .S(_1226__bF_buf0) );
MU2IX1 MU2IX1_92 ( .gnd!(gnd!), .vdd!(vdd!), .IN0(_849_), .IN1(_844_), .Q(_850_), .S(_1221__bF_buf0) );
ON21X1 ON21X1_260 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1576_), .B(_1221__bF_buf1), .C(_2034_), .Q(_851_) );
AN21X1 AN21X1_135 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1579_), .B(_1941_), .C(_866__bF_buf1), .Q(_852_) );
AN22X1 AN22X1_47 ( .gnd!(gnd!), .vdd!(vdd!), .A(_852_), .B(_851_), .C(_866__bF_buf1), .D(_850_), .Q(_853_) );
ON211X1 ON211X1_70 ( .gnd!(gnd!), .vdd!(vdd!), .A(_952__bF_buf0), .B(_853_), .C(_843_), .D(_909__bF_buf3), .Q(_854_) );
AN22X1 AN22X1_48 ( .gnd!(gnd!), .vdd!(vdd!), .A(_866__bF_buf0), .B(_1524__bF_buf0), .C(_854_), .D(_824_), .Q(ALU_r_22_) );
AN22X1 AN22X1_49 ( .gnd!(gnd!), .vdd!(vdd!), .A(_804_), .B(_827_), .C(_764_), .D(_825_), .Q(_857_) );
NA2X1 NA2X1_468 ( .gnd!(gnd!), .vdd!(vdd!), .A(_837_), .B(_836_), .Q(_858_) );
NO2X1 NO2X1_179 ( .gnd!(gnd!), .vdd!(vdd!), .A(_835_), .B(_858_), .Q(_859_) );
INX1 INX1_129 ( .gnd!(gnd!), .vdd!(vdd!), .A(_859_), .Q(_860_) );
INX1 INX1_130 ( .gnd!(gnd!), .vdd!(vdd!), .A(_841_), .Q(_861_) );
INX1 INX1_131 ( .gnd!(gnd!), .vdd!(vdd!), .A(ALU_a_23_), .Q(_862_) );
NA2X1 NA2X1_469 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1212__bF_buf2), .B(ALU_b_23_), .Q(_863_) );
INX1 INX1_132 ( .gnd!(gnd!), .vdd!(vdd!), .A(ALU_b_23_), .Q(_864_) );
NA2X1 NA2X1_470 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1059__bF_buf2), .B(_864_), .Q(_865_) );
NA2X1 NA2X1_471 ( .gnd!(gnd!), .vdd!(vdd!), .A(_865_), .B(_863_), .Q(_867_) );
NO2X1 NO2X1_180 ( .gnd!(gnd!), .vdd!(vdd!), .A(_862_), .B(_867_), .Q(_868_) );
NA2X1 NA2X1_472 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1212__bF_buf2), .B(_864_), .Q(_869_) );
NA2X1 NA2X1_473 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1059__bF_buf2), .B(ALU_b_23_), .Q(_870_) );
NA3I1X1 NA3I1X1_90 ( .gnd!(gnd!), .vdd!(vdd!), .AN(ALU_a_23_), .B(_869_), .C(_870_), .Q(_871_) );
INX1 INX1_133 ( .gnd!(gnd!), .vdd!(vdd!), .A(_871_), .Q(_872_) );
ON221X1 ON221X1_2 ( .gnd!(gnd!), .vdd!(vdd!), .A(_868_), .B(_872_), .C(_861_), .D(_857_), .E(_860_), .Q(_873_) );
NA3I1X1 NA3I1X1_91 ( .gnd!(gnd!), .vdd!(vdd!), .AN(_862_), .B(_863_), .C(_865_), .Q(_874_) );
ON211X1 ON211X1_71 ( .gnd!(gnd!), .vdd!(vdd!), .A(_840_), .B(_859_), .C(_874_), .D(_871_), .Q(_875_) );
NA3I1X1 NA3I1X1_92 ( .gnd!(gnd!), .vdd!(vdd!), .AN(_941__bF_buf1), .B(_873_), .C(_875_), .Q(_876_) );
NO2X1 NO2X1_181 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1227__bF_buf5), .B(_1947_), .Q(_878_) );
MU2IX1 MU2IX1_93 ( .gnd!(gnd!), .vdd!(vdd!), .IN0(ALU_a_23_), .IN1(ALU_a_22_), .Q(_879_), .S(_1235__bF_buf1) );
MU2X1 MU2X1_199 ( .gnd!(gnd!), .vdd!(vdd!), .IN0(_810_), .IN1(_879_), .Q(_880_), .S(_1233__bF_buf3) );
NA2X1 NA2X1_474 ( .gnd!(gnd!), .vdd!(vdd!), .A(_880_), .B(_1252__bF_buf0), .Q(_881_) );
ON21X1 ON21X1_261 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1252__bF_buf0), .B(_744_), .C(_881_), .Q(_882_) );
NA2X1 NA2X1_475 ( .gnd!(gnd!), .vdd!(vdd!), .A(_882_), .B(_1227__bF_buf0), .Q(_883_) );
NA2X1 NA2X1_476 ( .gnd!(gnd!), .vdd!(vdd!), .A(_883_), .B(_1222__bF_buf3), .Q(_884_) );
ON22X1 ON22X1_40 ( .gnd!(gnd!), .vdd!(vdd!), .A(_884_), .B(_878_), .C(_1222__bF_buf2), .D(_1653_), .Q(_885_) );
NA2X1 NA2X1_477 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1642_), .B(_1222__bF_buf1), .Q(_886_) );
NA2X1 NA2X1_478 ( .gnd!(gnd!), .vdd!(vdd!), .A(_886_), .B(_2034_), .Q(_887_) );
NA2X1 NA2X1_479 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1639_), .B(_712_), .Q(_889_) );
AN31X1 AN31X1_55 ( .gnd!(gnd!), .vdd!(vdd!), .A(EXT_type_bF_buf1), .B(_889_), .C(_887_), .D(_952__bF_buf0), .Q(_890_) );
ON21X1 ON21X1_262 ( .gnd!(gnd!), .vdd!(vdd!), .A(EXT_type_bF_buf2), .B(_885_), .C(_890_), .Q(_891_) );
AN21X1 AN21X1_136 ( .gnd!(gnd!), .vdd!(vdd!), .A(_862_), .B(_864_), .C(_1330_), .Q(_892_) );
ON31X1 ON31X1_45 ( .gnd!(gnd!), .vdd!(vdd!), .A(_862_), .B(_864_), .C(_1328__bF_buf0), .D(_892_), .Q(_893_) );
ON31X1 ON31X1_46 ( .gnd!(gnd!), .vdd!(vdd!), .A(_862_), .B(_864_), .C(_1526__bF_buf3), .D(_893_), .Q(_894_) );
ON21X1 ON21X1_263 ( .gnd!(gnd!), .vdd!(vdd!), .A(_894_), .B(_909__bF_buf0), .C(_1143__bF_buf1), .Q(_895_) );
AN31X1 AN31X1_56 ( .gnd!(gnd!), .vdd!(vdd!), .A(_909__bF_buf1), .B(_876_), .C(_891_), .D(_895_), .Q(ALU_r_23_) );
NA2X1 NA2X1_480 ( .gnd!(gnd!), .vdd!(vdd!), .A(ALU_a_24_), .B(ALU_b_24_), .Q(_896_) );
NO2X1 NO2X1_182 ( .gnd!(gnd!), .vdd!(vdd!), .A(_896_), .B(_1328__bF_buf2), .Q(_897_) );
ON22X1 ON22X1_41 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1329__bF_buf3), .B(_888__bF_buf0), .C(ALU_a_24_), .D(ALU_b_24_), .Q(_899_) );
ON22X1 ON22X1_42 ( .gnd!(gnd!), .vdd!(vdd!), .A(_897_), .B(_899_), .C(_1526__bF_buf4), .D(_896_), .Q(_900_) );
NA2X1 NA2X1_481 ( .gnd!(gnd!), .vdd!(vdd!), .A(_900_), .B(_1525__bF_buf4), .Q(_901_) );
AN21X1 AN21X1_137 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1222__bF_buf4), .B(_1695_), .C(_2033_), .Q(_902_) );
NO2I1X1 NO2I1X1_36 ( .gnd!(gnd!), .vdd!(vdd!), .AN(_1694_), .B(_902_), .Q(_903_) );
AND2X2 AND2X2_31 ( .gnd!(gnd!), .vdd!(vdd!), .A(_776_), .B(_1230__bF_buf0), .Q(_904_) );
NA2X1 NA2X1_482 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1334_), .B(_1338_), .Q(_905_) );
MU2X1 MU2X1_200 ( .gnd!(gnd!), .vdd!(vdd!), .IN0(_905_), .IN1(_845_), .Q(_906_), .S(_1240__bF_buf2) );
ON21X1 ON21X1_264 ( .gnd!(gnd!), .vdd!(vdd!), .A(_906_), .B(_1230__bF_buf0), .C(_1227__bF_buf0), .Q(_907_) );
ON22X1 ON22X1_43 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1964_), .B(_1227__bF_buf0), .C(_904_), .D(_907_), .Q(_908_) );
MU2IX1 MU2IX1_94 ( .gnd!(gnd!), .vdd!(vdd!), .IN0(_1688_), .IN1(_908_), .Q(_910_), .S(_1222__bF_buf0) );
ON22X1 ON22X1_44 ( .gnd!(gnd!), .vdd!(vdd!), .A(_910_), .B(EXT_type_bF_buf6), .C(_1942_), .D(_903_), .Q(_911_) );
ON211X1 ON211X1_72 ( .gnd!(gnd!), .vdd!(vdd!), .A(_838_), .B(_832_), .C(_874_), .D(_871_), .Q(_912_) );
NA2I1X1 NA2I1X1_55 ( .gnd!(gnd!), .vdd!(vdd!), .AN(_912_), .B(_825_), .Q(_913_) );
NO2X1 NO2X1_183 ( .gnd!(gnd!), .vdd!(vdd!), .A(_913_), .B(_763_), .Q(_914_) );
ON21X1 ON21X1_265 ( .gnd!(gnd!), .vdd!(vdd!), .A(_859_), .B(_868_), .C(_871_), .Q(_915_) );
ON221X1 ON221X1_3 ( .gnd!(gnd!), .vdd!(vdd!), .A(_828_), .B(_912_), .C(_913_), .D(_762_), .E(_915_), .Q(_916_) );
AN21X1 AN21X1_138 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1983_), .B(_914_), .C(_916_), .Q(_917_) );
EN2X1 EN2X1_1 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1059__bF_buf3), .B(ALU_b_24_), .Q(_918_) );
NA2I1X1 NA2I1X1_56 ( .gnd!(gnd!), .vdd!(vdd!), .AN(ALU_a_24_), .B(_918_), .Q(_919_) );
NA2I1X1 NA2I1X1_57 ( .gnd!(gnd!), .vdd!(vdd!), .AN(_918_), .B(ALU_a_24_), .Q(_921_) );
AND2X2 AND2X2_32 ( .gnd!(gnd!), .vdd!(vdd!), .A(_921_), .B(_919_), .Q(_922_) );
NA2X1 NA2X1_483 ( .gnd!(gnd!), .vdd!(vdd!), .A(_917_), .B(_922_), .Q(_923_) );
NO3X1 NO3X1_5 ( .gnd!(gnd!), .vdd!(vdd!), .A(_912_), .B(_771_), .C(_805_), .Q(_924_) );
NA2X1 NA2X1_484 ( .gnd!(gnd!), .vdd!(vdd!), .A(_793_), .B(_924_), .Q(_925_) );
NA2X1 NA2X1_485 ( .gnd!(gnd!), .vdd!(vdd!), .A(_760_), .B(_737_), .Q(_926_) );
ON31X1 ON31X1_47 ( .gnd!(gnd!), .vdd!(vdd!), .A(_701_), .B(_740_), .C(_696_), .D(_926_), .Q(_927_) );
ON21X1 ON21X1_266 ( .gnd!(gnd!), .vdd!(vdd!), .A(_912_), .B(_828_), .C(_915_), .Q(_928_) );
AN21X1 AN21X1_139 ( .gnd!(gnd!), .vdd!(vdd!), .A(_927_), .B(_924_), .C(_928_), .Q(_929_) );
ON21X1 ON21X1_267 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2001_), .B(_925_), .C(_929_), .Q(_930_) );
NA2X1 NA2X1_486 ( .gnd!(gnd!), .vdd!(vdd!), .A(_921_), .B(_919_), .Q(_932_) );
NA2X1 NA2X1_487 ( .gnd!(gnd!), .vdd!(vdd!), .A(_930_), .B(_932_), .Q(_933_) );
NA2X1 NA2X1_488 ( .gnd!(gnd!), .vdd!(vdd!), .A(_923_), .B(_933_), .Q(_934_) );
NA2X1 NA2X1_489 ( .gnd!(gnd!), .vdd!(vdd!), .A(_934_), .B(_952__bF_buf3), .Q(_935_) );
ON211X1 ON211X1_73 ( .gnd!(gnd!), .vdd!(vdd!), .A(_952__bF_buf5), .B(_911_), .C(_935_), .D(_909__bF_buf3), .Q(_936_) );
AN22X1 AN22X1_50 ( .gnd!(gnd!), .vdd!(vdd!), .A(_866__bF_buf3), .B(_1524__bF_buf2), .C(_936_), .D(_901_), .Q(ALU_r_24_) );
NA2X1 NA2X1_490 ( .gnd!(gnd!), .vdd!(vdd!), .A(ALU_a_25_), .B(ALU_b_25_), .Q(_937_) );
NO2X1 NO2X1_184 ( .gnd!(gnd!), .vdd!(vdd!), .A(_937_), .B(_1328__bF_buf2), .Q(_938_) );
ON22X1 ON22X1_45 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1329__bF_buf1), .B(_888__bF_buf0), .C(ALU_a_25_), .D(ALU_b_25_), .Q(_939_) );
ON22X1 ON22X1_46 ( .gnd!(gnd!), .vdd!(vdd!), .A(_938_), .B(_939_), .C(_1526__bF_buf4), .D(_937_), .Q(_940_) );
NA2X1 NA2X1_491 ( .gnd!(gnd!), .vdd!(vdd!), .A(_940_), .B(_1525__bF_buf1), .Q(_942_) );
NA2X1 NA2X1_492 ( .gnd!(gnd!), .vdd!(vdd!), .A(_918_), .B(ALU_a_24_), .Q(_943_) );
EN2X1 EN2X1_2 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1212__bF_buf3), .B(ALU_b_25_), .Q(_944_) );
NA2I1X1 NA2I1X1_58 ( .gnd!(gnd!), .vdd!(vdd!), .AN(_944_), .B(ALU_a_25_), .Q(_945_) );
NA2I1X1 NA2I1X1_59 ( .gnd!(gnd!), .vdd!(vdd!), .AN(ALU_a_25_), .B(_944_), .Q(_946_) );
NA2X1 NA2X1_493 ( .gnd!(gnd!), .vdd!(vdd!), .A(_945_), .B(_946_), .Q(_947_) );
NA3I1X1 NA3I1X1_93 ( .gnd!(gnd!), .vdd!(vdd!), .AN(_947_), .B(_943_), .C(_933_), .Q(_948_) );
INX1 INX1_134 ( .gnd!(gnd!), .vdd!(vdd!), .A(_943_), .Q(_949_) );
NA2X1 NA2X1_494 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1983_), .B(_914_), .Q(_950_) );
AN22X1 AN22X1_51 ( .gnd!(gnd!), .vdd!(vdd!), .A(_919_), .B(_921_), .C(_950_), .D(_929_), .Q(_951_) );
ON21X1 ON21X1_268 ( .gnd!(gnd!), .vdd!(vdd!), .A(_951_), .B(_949_), .C(_947_), .Q(_953_) );
NO3X1 NO3X1_6 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1269_), .B(_1226__bF_buf1), .C(_2036_), .Q(_954_) );
NO2X1 NO2X1_185 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2033_), .B(_1705_), .Q(_955_) );
ON31X1 ON31X1_48 ( .gnd!(gnd!), .vdd!(vdd!), .A(_902_), .B(_954_), .C(_955_), .D(EXT_type_bF_buf4), .Q(_956_) );
MU2IX1 MU2IX1_95 ( .gnd!(gnd!), .vdd!(vdd!), .IN0(ALU_a_25_), .IN1(ALU_a_24_), .Q(_957_), .S(_1235__bF_buf4) );
MU2IX1 MU2IX1_96 ( .gnd!(gnd!), .vdd!(vdd!), .IN0(_879_), .IN1(_957_), .Q(_958_), .S(_1233__bF_buf3) );
MU2IX1 MU2IX1_97 ( .gnd!(gnd!), .vdd!(vdd!), .IN0(_811_), .IN1(_958_), .Q(_959_), .S(_1252__bF_buf0) );
MU2IX1 MU2IX1_98 ( .gnd!(gnd!), .vdd!(vdd!), .IN0(_959_), .IN1(_2028_), .Q(_960_), .S(_1226__bF_buf0) );
NA2X1 NA2X1_495 ( .gnd!(gnd!), .vdd!(vdd!), .A(_960_), .B(_1322__bF_buf3), .Q(_961_) );
ON311X1 ON311X1_5 ( .gnd!(gnd!), .vdd!(vdd!), .A(EXT_type_bF_buf2), .B(_1222__bF_buf3), .C(_1715_), .D(_961_), .E(_956_), .Q(_962_) );
NO2X1 NO2X1_186 ( .gnd!(gnd!), .vdd!(vdd!), .A(_952__bF_buf2), .B(_962_), .Q(_964_) );
AO311X1 AO311X1_2 ( .gnd!(gnd!), .vdd!(vdd!), .A(_952__bF_buf2), .B(_948_), .C(_953_), .D(_1525__bF_buf2), .E(_964_), .Q(_965_) );
AN22X1 AN22X1_52 ( .gnd!(gnd!), .vdd!(vdd!), .A(_866__bF_buf2), .B(_1524__bF_buf3), .C(_965_), .D(_942_), .Q(ALU_r_25_) );
NA2X1 NA2X1_496 ( .gnd!(gnd!), .vdd!(vdd!), .A(ALU_a_26_), .B(ALU_b_26_), .Q(_966_) );
NO2X1 NO2X1_187 ( .gnd!(gnd!), .vdd!(vdd!), .A(_966_), .B(_1328__bF_buf2), .Q(_967_) );
ON22X1 ON22X1_47 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1329__bF_buf1), .B(_888__bF_buf0), .C(ALU_a_26_), .D(ALU_b_26_), .Q(_968_) );
ON22X1 ON22X1_48 ( .gnd!(gnd!), .vdd!(vdd!), .A(_967_), .B(_968_), .C(_1526__bF_buf3), .D(_966_), .Q(_969_) );
NA2X1 NA2X1_497 ( .gnd!(gnd!), .vdd!(vdd!), .A(_969_), .B(_1525__bF_buf3), .Q(_970_) );
EN2X1 EN2X1_3 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1212__bF_buf1), .B(ALU_b_26_), .Q(_971_) );
NA2I1X1 NA2I1X1_60 ( .gnd!(gnd!), .vdd!(vdd!), .AN(_971_), .B(ALU_a_26_), .Q(_972_) );
NA2I1X1 NA2I1X1_61 ( .gnd!(gnd!), .vdd!(vdd!), .AN(ALU_a_26_), .B(_971_), .Q(_974_) );
NA2X1 NA2X1_498 ( .gnd!(gnd!), .vdd!(vdd!), .A(_972_), .B(_974_), .Q(_975_) );
NO2X1 NO2X1_188 ( .gnd!(gnd!), .vdd!(vdd!), .A(_947_), .B(_922_), .Q(_976_) );
NA2X1 NA2X1_499 ( .gnd!(gnd!), .vdd!(vdd!), .A(_930_), .B(_976_), .Q(_977_) );
NA2X1 NA2X1_500 ( .gnd!(gnd!), .vdd!(vdd!), .A(_945_), .B(_943_), .Q(_978_) );
NA2X1 NA2X1_501 ( .gnd!(gnd!), .vdd!(vdd!), .A(_978_), .B(_946_), .Q(_979_) );
AN21X1 AN21X1_140 ( .gnd!(gnd!), .vdd!(vdd!), .A(_977_), .B(_979_), .C(_975_), .Q(_980_) );
EN2X1 EN2X1_4 ( .gnd!(gnd!), .vdd!(vdd!), .A(_971_), .B(ALU_a_26_), .Q(_981_) );
NA2I1X1 NA2I1X1_62 ( .gnd!(gnd!), .vdd!(vdd!), .AN(_947_), .B(_932_), .Q(_982_) );
ON21X1 ON21X1_269 ( .gnd!(gnd!), .vdd!(vdd!), .A(_917_), .B(_982_), .C(_979_), .Q(_983_) );
NO2X1 NO2X1_189 ( .gnd!(gnd!), .vdd!(vdd!), .A(_981_), .B(_983_), .Q(_985_) );
ON21X1 ON21X1_270 ( .gnd!(gnd!), .vdd!(vdd!), .A(_985_), .B(_980_), .C(_952__bF_buf3), .Q(_986_) );
AND2X2 AND2X2_33 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1742_), .B(_1960_), .Q(_987_) );
NO2X1 NO2X1_190 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2033_), .B(_1745_), .Q(_988_) );
NO2X1 NO2X1_191 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2036_), .B(_1743_), .Q(_989_) );
ON31X1 ON31X1_49 ( .gnd!(gnd!), .vdd!(vdd!), .A(_902_), .B(_989_), .C(_988_), .D(EXT_type_bF_buf1), .Q(_990_) );
NA2X1 NA2X1_502 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1353_), .B(_1335_), .Q(_991_) );
MU2IX1 MU2IX1_99 ( .gnd!(gnd!), .vdd!(vdd!), .IN0(_991_), .IN1(_905_), .Q(_992_), .S(_1240__bF_buf2) );
AND2X2 AND2X2_34 ( .gnd!(gnd!), .vdd!(vdd!), .A(_992_), .B(_1252__bF_buf3), .Q(_993_) );
ON21X1 ON21X1_271 ( .gnd!(gnd!), .vdd!(vdd!), .A(_846_), .B(_1252__bF_buf0), .C(_1227__bF_buf0), .Q(_994_) );
ON22X1 ON22X1_49 ( .gnd!(gnd!), .vdd!(vdd!), .A(_706_), .B(_1227__bF_buf0), .C(_994_), .D(_993_), .Q(_996_) );
NA2X1 NA2X1_503 ( .gnd!(gnd!), .vdd!(vdd!), .A(_996_), .B(_1322__bF_buf0), .Q(_997_) );
NA2X1 NA2X1_504 ( .gnd!(gnd!), .vdd!(vdd!), .A(_990_), .B(_997_), .Q(_998_) );
ON311X1 ON311X1_6 ( .gnd!(gnd!), .vdd!(vdd!), .A(_952__bF_buf5), .B(_987_), .C(_998_), .D(_909__bF_buf3), .E(_986_), .Q(_999_) );
AN22X1 AN22X1_53 ( .gnd!(gnd!), .vdd!(vdd!), .A(_866__bF_buf0), .B(_1524__bF_buf0), .C(_999_), .D(_970_), .Q(ALU_r_26_) );
NA2X1 NA2X1_505 ( .gnd!(gnd!), .vdd!(vdd!), .A(ALU_a_27_), .B(ALU_b_27_), .Q(_1000_) );
NO2X1 NO2X1_192 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1000_), .B(_1328__bF_buf1), .Q(_1001_) );
ON22X1 ON22X1_50 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1329__bF_buf0), .B(_888__bF_buf3), .C(ALU_a_27_), .D(ALU_b_27_), .Q(_1002_) );
ON22X1 ON22X1_51 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1001_), .B(_1002_), .C(_1526__bF_buf4), .D(_1000_), .Q(_1003_) );
NA2X1 NA2X1_506 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1003_), .B(_1525__bF_buf1), .Q(_1004_) );
NA2X1 NA2X1_507 ( .gnd!(gnd!), .vdd!(vdd!), .A(_983_), .B(_981_), .Q(_1006_) );
NA2X1 NA2X1_508 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1006_), .B(_972_), .Q(_1007_) );
EN2X1 EN2X1_5 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1059__bF_buf3), .B(ALU_b_27_), .Q(_1008_) );
NA2X1 NA2X1_509 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1008_), .B(ALU_a_27_), .Q(_1009_) );
EN2X1 EN2X1_6 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1212__bF_buf1), .B(ALU_b_27_), .Q(_1010_) );
NA2I1X1 NA2I1X1_63 ( .gnd!(gnd!), .vdd!(vdd!), .AN(ALU_a_27_), .B(_1010_), .Q(_1011_) );
NA2X1 NA2X1_510 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1009_), .B(_1011_), .Q(_1012_) );
NO2X1 NO2X1_193 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1012_), .B(_1007_), .Q(_1013_) );
AN22X1 AN22X1_54 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1009_), .B(_1011_), .C(_1006_), .D(_972_), .Q(_1014_) );
NO2X1 NO2X1_194 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2036_), .B(_1778_), .Q(_1015_) );
NO2X1 NO2X1_195 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2033_), .B(_1776_), .Q(_1017_) );
ON31X1 ON31X1_50 ( .gnd!(gnd!), .vdd!(vdd!), .A(_902_), .B(_1017_), .C(_1015_), .D(EXT_type_bF_buf4), .Q(_1018_) );
NA2X1 NA2X1_511 ( .gnd!(gnd!), .vdd!(vdd!), .A(_745_), .B(_1226__bF_buf0), .Q(_1019_) );
NA2X1 NA2X1_512 ( .gnd!(gnd!), .vdd!(vdd!), .A(_957_), .B(_1240__bF_buf2), .Q(_1020_) );
MU2X1 MU2X1_201 ( .gnd!(gnd!), .vdd!(vdd!), .IN0(ALU_a_27_), .IN1(ALU_a_26_), .Q(_1021_), .S(_1235__bF_buf4) );
ON21X1 ON21X1_272 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1240__bF_buf2), .B(_1021_), .C(_1020_), .Q(_1022_) );
MU2IX1 MU2IX1_100 ( .gnd!(gnd!), .vdd!(vdd!), .IN0(_880_), .IN1(_1022_), .Q(_1023_), .S(_1252__bF_buf0) );
ON211X1 ON211X1_74 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1226__bF_buf0), .B(_1023_), .C(_1019_), .D(_1322__bF_buf3), .Q(_1024_) );
AN21X1 AN21X1_141 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1787_), .B(_1960_), .C(_952__bF_buf0), .Q(_1025_) );
AN31X1 AN31X1_57 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1024_), .B(_1025_), .C(_1018_), .D(_1525__bF_buf2), .Q(_1026_) );
ON31X1 ON31X1_51 ( .gnd!(gnd!), .vdd!(vdd!), .A(_941__bF_buf1), .B(_1014_), .C(_1013_), .D(_1026_), .Q(_1028_) );
AN22X1 AN22X1_55 ( .gnd!(gnd!), .vdd!(vdd!), .A(_866__bF_buf3), .B(_1524__bF_buf2), .C(_1028_), .D(_1004_), .Q(ALU_r_27_) );
NA2X1 NA2X1_513 ( .gnd!(gnd!), .vdd!(vdd!), .A(ALU_a_28_), .B(ALU_b_28_), .Q(_1029_) );
NO2X1 NO2X1_196 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1029_), .B(_1328__bF_buf2), .Q(_1030_) );
ON22X1 ON22X1_52 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1329__bF_buf1), .B(_888__bF_buf0), .C(ALU_a_28_), .D(ALU_b_28_), .Q(_1031_) );
ON22X1 ON22X1_53 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1030_), .B(_1031_), .C(_1526__bF_buf4), .D(_1029_), .Q(_1032_) );
NA2X1 NA2X1_514 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1032_), .B(_1525__bF_buf1), .Q(_1033_) );
NO2X1 NO2X1_197 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1012_), .B(_975_), .Q(_1034_) );
NA2X1 NA2X1_515 ( .gnd!(gnd!), .vdd!(vdd!), .A(_976_), .B(_1034_), .Q(_1035_) );
NA2X1 NA2X1_516 ( .gnd!(gnd!), .vdd!(vdd!), .A(_972_), .B(_1009_), .Q(_1036_) );
AN32X1 AN32X1_4 ( .gnd!(gnd!), .vdd!(vdd!), .A(_946_), .B(_978_), .C(_1034_), .D(_1011_), .E(_1036_), .Q(_1038_) );
ON21X1 ON21X1_273 ( .gnd!(gnd!), .vdd!(vdd!), .A(_917_), .B(_1035_), .C(_1038_), .Q(_1039_) );
EN2X1 EN2X1_7 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1212__bF_buf3), .B(ALU_b_28_), .Q(_1040_) );
NA2I1X1 NA2I1X1_64 ( .gnd!(gnd!), .vdd!(vdd!), .AN(_1040_), .B(ALU_a_28_), .Q(_1041_) );
NA2I1X1 NA2I1X1_65 ( .gnd!(gnd!), .vdd!(vdd!), .AN(ALU_a_28_), .B(_1040_), .Q(_1042_) );
NA2X1 NA2X1_517 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1041_), .B(_1042_), .Q(_1043_) );
NA2X1 NA2X1_518 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1039_), .B(_1043_), .Q(_1044_) );
AND2X2 AND2X2_35 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1009_), .B(_1011_), .Q(_1045_) );
NA2X1 NA2X1_519 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1045_), .B(_981_), .Q(_1046_) );
NO2X1 NO2X1_198 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1046_), .B(_982_), .Q(_1047_) );
ON221X1 ON221X1_4 ( .gnd!(gnd!), .vdd!(vdd!), .A(_972_), .B(_1012_), .C(_979_), .D(_1046_), .E(_1009_), .Q(_1049_) );
AN21X1 AN21X1_142 ( .gnd!(gnd!), .vdd!(vdd!), .A(_930_), .B(_1047_), .C(_1049_), .Q(_1050_) );
INX1 INX1_135 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1043_), .Q(_1051_) );
NA2X1 NA2X1_520 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1050_), .B(_1051_), .Q(_1052_) );
NA2X1 NA2X1_521 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1044_), .B(_1052_), .Q(_1053_) );
AND3X4 AND3X4_6 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1832_), .B(_1222__bF_buf1), .C(_1833_), .Q(_1054_) );
ON22X1 ON22X1_54 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1054_), .B(_2033_), .C(_1832_), .D(_2036_), .Q(_1055_) );
AND2X2 AND2X2_36 ( .gnd!(gnd!), .vdd!(vdd!), .A(_777_), .B(_1226__bF_buf0), .Q(_1056_) );
NA2I1X1 NA2I1X1_66 ( .gnd!(gnd!), .vdd!(vdd!), .AN(_991_), .B(_1240__bF_buf2), .Q(_1057_) );
AN31X1 AN31X1_58 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1354_), .B(_1349_), .C(_1233__bF_buf1), .D(_1230__bF_buf0), .Q(_1058_) );
AN22X1 AN22X1_56 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1057_), .B(_1058_), .C(_906_), .D(_1230__bF_buf0), .Q(_1060_) );
AN211X1 AN211X1_8 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1227__bF_buf6), .B(_1060_), .C(_1400_), .D(_1056_), .Q(_1061_) );
AN221X1 AN221X1_7 ( .gnd!(gnd!), .vdd!(vdd!), .A(EXT_type_bF_buf6), .B(_1055_), .C(_1840_), .D(_1960_), .E(_1061_), .Q(_1062_) );
NA2X1 NA2X1_522 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1062_), .B(_941__bF_buf4), .Q(_1063_) );
ON211X1 ON211X1_75 ( .gnd!(gnd!), .vdd!(vdd!), .A(_941__bF_buf1), .B(_1053_), .C(_1063_), .D(_909__bF_buf4), .Q(_1064_) );
AN22X1 AN22X1_57 ( .gnd!(gnd!), .vdd!(vdd!), .A(_866__bF_buf2), .B(_1524__bF_buf3), .C(_1064_), .D(_1033_), .Q(ALU_r_28_) );
NA2X1 NA2X1_523 ( .gnd!(gnd!), .vdd!(vdd!), .A(ALU_a_29_), .B(ALU_b_29_), .Q(_1065_) );
NO2X1 NO2X1_199 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1065_), .B(_1328__bF_buf2), .Q(_1066_) );
ON22X1 ON22X1_55 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1329__bF_buf1), .B(_888__bF_buf4), .C(ALU_a_29_), .D(ALU_b_29_), .Q(_1067_) );
ON22X1 ON22X1_56 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1066_), .B(_1067_), .C(_1526__bF_buf3), .D(_1065_), .Q(_1068_) );
NA2X1 NA2X1_524 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1068_), .B(_1525__bF_buf4), .Q(_1070_) );
EN2X1 EN2X1_8 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1212__bF_buf3), .B(ALU_b_29_), .Q(_1071_) );
NA2I1X1 NA2I1X1_67 ( .gnd!(gnd!), .vdd!(vdd!), .AN(_1071_), .B(ALU_a_29_), .Q(_1072_) );
NA2I1X1 NA2I1X1_68 ( .gnd!(gnd!), .vdd!(vdd!), .AN(ALU_a_29_), .B(_1071_), .Q(_1073_) );
NA2X1 NA2X1_525 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1072_), .B(_1073_), .Q(_1074_) );
ON211X1 ON211X1_76 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1050_), .B(_1043_), .C(_1041_), .D(_1074_), .Q(_1075_) );
ON21X1 ON21X1_274 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1050_), .B(_1043_), .C(_1041_), .Q(_1076_) );
INX1 INX1_136 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1074_), .Q(_1077_) );
NA2X1 NA2X1_526 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1076_), .B(_1077_), .Q(_1078_) );
NO2X1 NO2X1_200 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1221__bF_buf2), .B(_1862_), .Q(_1079_) );
NO2X1 NO2X1_201 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2033_), .B(_1079_), .Q(_1081_) );
NO2X1 NO2X1_202 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2036_), .B(_1863_), .Q(_1082_) );
ON21X1 ON21X1_275 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1081_), .B(_1082_), .C(EXT_type_bF_buf4), .Q(_1083_) );
NA2X1 NA2X1_527 ( .gnd!(gnd!), .vdd!(vdd!), .A(_812_), .B(_1226__bF_buf6), .Q(_1084_) );
NA2I1X1 NA2I1X1_69 ( .gnd!(gnd!), .vdd!(vdd!), .AN(_1021_), .B(_1240__bF_buf2), .Q(_1085_) );
MU2IX1 MU2IX1_101 ( .gnd!(gnd!), .vdd!(vdd!), .IN0(ALU_a_29_), .IN1(ALU_a_28_), .Q(_1086_), .S(_1235__bF_buf4) );
AN21X1 AN21X1_143 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1086_), .B(_1233__bF_buf3), .C(_1230__bF_buf1), .Q(_1087_) );
AO22X2 AO22X2_28 ( .gnd!(gnd!), .vdd!(vdd!), .A(_958_), .B(_1230__bF_buf1), .C(_1085_), .D(_1087_), .Q(_1088_) );
ON211X1 ON211X1_77 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1226__bF_buf0), .B(_1088_), .C(_1084_), .D(_1322__bF_buf3), .Q(_1089_) );
NA2X1 NA2X1_528 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1873_), .B(_1960_), .Q(_1090_) );
AN31X1 AN31X1_59 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1089_), .B(_1090_), .C(_1083_), .D(_952__bF_buf0), .Q(_1092_) );
AN31X1 AN31X1_60 ( .gnd!(gnd!), .vdd!(vdd!), .A(_952__bF_buf2), .B(_1075_), .C(_1078_), .D(_1092_), .Q(_1093_) );
NA2I1X1 NA2I1X1_70 ( .gnd!(gnd!), .vdd!(vdd!), .AN(_1093_), .B(_909__bF_buf1), .Q(_1094_) );
AN22X1 AN22X1_58 ( .gnd!(gnd!), .vdd!(vdd!), .A(_866__bF_buf5), .B(_1524__bF_buf1), .C(_1094_), .D(_1070_), .Q(ALU_r_29_) );
NA2X1 NA2X1_529 ( .gnd!(gnd!), .vdd!(vdd!), .A(ALU_a_30_), .B(ALU_b_30_), .Q(_1095_) );
NO2X1 NO2X1_203 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1095_), .B(_1328__bF_buf2), .Q(_1096_) );
ON22X1 ON22X1_57 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1329__bF_buf3), .B(_888__bF_buf0), .C(ALU_a_30_), .D(ALU_b_30_), .Q(_1097_) );
ON22X1 ON22X1_58 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1096_), .B(_1097_), .C(_1526__bF_buf4), .D(_1095_), .Q(_1098_) );
NA2X1 NA2X1_530 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1098_), .B(_1525__bF_buf4), .Q(_1099_) );
NO2X1 NO2X1_204 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1043_), .B(_1074_), .Q(_1100_) );
INX1 INX1_137 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1100_), .Q(_1102_) );
ON21X1 ON21X1_276 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1074_), .B(_1041_), .C(_1072_), .Q(_1103_) );
INX1 INX1_138 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1103_), .Q(_1104_) );
ON21X1 ON21X1_277 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1050_), .B(_1102_), .C(_1104_), .Q(_1105_) );
EN2X1 EN2X1_9 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1212__bF_buf3), .B(ALU_b_30_), .Q(_1106_) );
NA2I1X1 NA2I1X1_71 ( .gnd!(gnd!), .vdd!(vdd!), .AN(_1106_), .B(ALU_a_30_), .Q(_1107_) );
NA2I1X1 NA2I1X1_72 ( .gnd!(gnd!), .vdd!(vdd!), .AN(ALU_a_30_), .B(_1106_), .Q(_1108_) );
NA2X1 NA2X1_531 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1107_), .B(_1108_), .Q(_1109_) );
INX1 INX1_139 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1109_), .Q(_1110_) );
NA2X1 NA2X1_532 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1105_), .B(_1110_), .Q(_1111_) );
AN21X1 AN21X1_144 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1039_), .B(_1100_), .C(_1103_), .Q(_1113_) );
NA2X1 NA2X1_533 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1113_), .B(_1109_), .Q(_1114_) );
NA2X1 NA2X1_534 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1114_), .B(_1111_), .Q(_1115_) );
NA2X1 NA2X1_535 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1115_), .B(_952__bF_buf5), .Q(_1116_) );
NO2X1 NO2X1_205 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1221__bF_buf1), .B(_1902_), .Q(_1117_) );
OA22X4 OA22X4_1 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1117_), .B(_2033_), .C(_1901_), .D(_2036_), .Q(_1118_) );
NA2X1 NA2X1_536 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1912_), .B(_1960_), .Q(_1119_) );
AND3X4 AND3X4_7 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1349_), .B(_1354_), .C(_1240__bF_buf5), .Q(_1120_) );
AO311X1 AO311X1_3 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1233__bF_buf1), .B(_1350_), .C(_1359_), .D(_1230__bF_buf0), .E(_1120_), .Q(_1121_) );
ON21X1 ON21X1_278 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1252__bF_buf3), .B(_992_), .C(_1121_), .Q(_1122_) );
MU2IX1 MU2IX1_102 ( .gnd!(gnd!), .vdd!(vdd!), .IN0(_1122_), .IN1(_848_), .Q(_1124_), .S(_1226__bF_buf0) );
OA221X1 OA221X1_1 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1400_), .B(_1124_), .C(_866__bF_buf4), .D(_1118_), .E(_1119_), .Q(_1125_) );
AN22X1 AN22X1_59 ( .gnd!(gnd!), .vdd!(vdd!), .A(_856_), .B(_898_), .C(_1125_), .D(_941__bF_buf2), .Q(_1126_) );
NA2X1 NA2X1_537 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1116_), .B(_1126_), .Q(_1127_) );
AN22X1 AN22X1_60 ( .gnd!(gnd!), .vdd!(vdd!), .A(_866__bF_buf3), .B(_1524__bF_buf2), .C(_1127_), .D(_1099_), .Q(ALU_r_30_) );
ON21X1 ON21X1_279 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1113_), .B(_1109_), .C(_1107_), .Q(_1128_) );
EN2X1 EN2X1_10 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1059__bF_buf2), .B(ALU_b_31_), .Q(_1129_) );
NA2X1 NA2X1_538 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1129_), .B(ALU_a_31_), .Q(_1130_) );
NA2I1X1 NA2I1X1_73 ( .gnd!(gnd!), .vdd!(vdd!), .AN(_1129_), .B(_1265_), .Q(_1131_) );
NA2X1 NA2X1_539 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1131_), .B(_1130_), .Q(_1132_) );
INX1 INX1_140 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1132_), .Q(_1134_) );
NA2X1 NA2X1_540 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1128_), .B(_1134_), .Q(_1135_) );
INX1 INX1_141 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1107_), .Q(_1136_) );
NA3I1X1 NA3I1X1_94 ( .gnd!(gnd!), .vdd!(vdd!), .AN(_1136_), .B(_1132_), .C(_1111_), .Q(_1137_) );
NA2X1 NA2X1_541 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1135_), .B(_1137_), .Q(_1138_) );
INX1 INX1_142 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1138_), .Q(ALU_sf) );
NA2X1 NA2X1_542 ( .gnd!(gnd!), .vdd!(vdd!), .A(ALU_a_31_), .B(ALU_b_31_), .Q(_1139_) );
NO2X1 NO2X1_206 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1139_), .B(_1328__bF_buf0), .Q(_1140_) );
ON22X1 ON22X1_59 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1329__bF_buf1), .B(_888__bF_buf4), .C(ALU_a_31_), .D(ALU_b_31_), .Q(_1141_) );
ON22X1 ON22X1_60 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1140_), .B(_1141_), .C(_1526__bF_buf3), .D(_1139_), .Q(_1142_) );
NA2X1 NA2X1_543 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1142_), .B(_1525__bF_buf0), .Q(_1144_) );
AN211X1 AN211X1_9 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1110_), .B(_1105_), .C(_1136_), .D(_1132_), .Q(_1145_) );
AN22X1 AN22X1_61 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1130_), .B(_1131_), .C(_1111_), .D(_1107_), .Q(_1146_) );
AND2X2 AND2X2_37 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1022_), .B(_1230__bF_buf0), .Q(_1147_) );
MU2IX1 MU2IX1_103 ( .gnd!(gnd!), .vdd!(vdd!), .IN0(_1086_), .IN1(_1257_), .Q(_1148_), .S(_1233__bF_buf3) );
ON31X1 ON31X1_52 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1230__bF_buf0), .B(_1437_), .C(_1148_), .D(_1227__bF_buf0), .Q(_1149_) );
ON22X1 ON22X1_61 ( .gnd!(gnd!), .vdd!(vdd!), .A(_882_), .B(_1227__bF_buf0), .C(_1147_), .D(_1149_), .Q(_1150_) );
AN31X1 AN31X1_61 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1227__bF_buf1), .B(_1637_), .C(_712_), .D(_1939_), .Q(_1151_) );
NO2X1 NO2X1_207 ( .gnd!(gnd!), .vdd!(vdd!), .A(_866__bF_buf1), .B(_1151_), .Q(_1152_) );
AN221X1 AN221X1_8 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1150_), .B(_1322__bF_buf1), .C(_1948_), .D(_1960_), .E(_1152_), .Q(_1153_) );
AN22X1 AN22X1_62 ( .gnd!(gnd!), .vdd!(vdd!), .A(_856_), .B(_898_), .C(_1153_), .D(_941__bF_buf2), .Q(_1155_) );
ON31X1 ON31X1_53 ( .gnd!(gnd!), .vdd!(vdd!), .A(_941__bF_buf0), .B(_1145_), .C(_1146_), .D(_1155_), .Q(_1156_) );
AN22X1 AN22X1_63 ( .gnd!(gnd!), .vdd!(vdd!), .A(_866__bF_buf5), .B(_1524__bF_buf1), .C(_1156_), .D(_1144_), .Q(ALU_r_31_) );
NA2X1 NA2X1_544 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1107_), .B(_1130_), .Q(_1157_) );
NA2X1 NA2X1_545 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1157_), .B(_1131_), .Q(_1158_) );
NA3I1X1 NA3I1X1_95 ( .gnd!(gnd!), .vdd!(vdd!), .AN(_1109_), .B(_1134_), .C(_1105_), .Q(_1159_) );
NA2X1 NA2X1_546 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1159_), .B(_1158_), .Q(ALU_cf) );
NO2X1 NO2X1_208 ( .gnd!(gnd!), .vdd!(vdd!), .A(ALU_a_0_), .B(ALU_b_0_), .Q(_1160_) );
NO2X1 NO2X1_209 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1160_), .B(_984_), .Q(_1161_) );
AN21X1 AN21X1_145 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1210_), .B(_1216_), .C(_1161_), .Q(_1162_) );
ON21X1 ON21X1_280 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1421_), .B(_1417_), .C(_1162_), .Q(_1164_) );
AN21X1 AN21X1_146 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1464_), .B(_1467_), .C(_1164_), .Q(_1165_) );
ON211X1 ON211X1_78 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1560_), .B(_1563_), .C(_1165_), .D(_1493_), .Q(_1166_) );
ON22X1 ON22X1_62 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1677_), .B(_1682_), .C(_1603_), .D(_1607_), .Q(_1167_) );
NO2X1 NO2X1_210 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1166_), .B(_1167_), .Q(_1168_) );
AN22X1 AN22X1_64 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1725_), .B(_1728_), .C(_1765_), .D(_1767_), .Q(_1169_) );
AND5X1 AND5X1_1 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1828_), .B(_1631_), .C(_2004_), .D(_1169_), .E(_1168_), .Q(_1170_) );
AN22X1 AN22X1_65 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2019_), .B(_2024_), .C(_1898_), .D(_1899_), .Q(_1171_) );
AN22X1 AN22X1_66 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1800_), .B(_1798_), .C(_1857_), .D(_1859_), .Q(_1172_) );
NA3X1 NA3X1_7 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1171_), .B(_1172_), .C(_1170_), .Q(_1173_) );
ON211X1 ON211X1_79 ( .gnd!(gnd!), .vdd!(vdd!), .A(_741_), .B(_739_), .C(_806_), .D(_807_), .Q(_1175_) );
AN22X1 AN22X1_67 ( .gnd!(gnd!), .vdd!(vdd!), .A(_700_), .B(_702_), .C(_773_), .D(_772_), .Q(_1176_) );
ON211X1 ON211X1_80 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1930_), .B(_1935_), .C(_1176_), .D(_934_), .Q(_1177_) );
NO3X1 NO3X1_7 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1177_), .B(_1173_), .C(_1175_), .Q(_1178_) );
NA3I1X1 NA3I1X1_96 ( .gnd!(gnd!), .vdd!(vdd!), .AN(_1045_), .B(_972_), .C(_1006_), .Q(_1179_) );
NA2X1 NA2X1_547 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1007_), .B(_1045_), .Q(_1180_) );
AN22X1 AN22X1_68 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1075_), .B(_1078_), .C(_1180_), .D(_1179_), .Q(_1181_) );
ON211X1 ON211X1_81 ( .gnd!(gnd!), .vdd!(vdd!), .A(_985_), .B(_980_), .C(_1044_), .D(_1052_), .Q(_1182_) );
ON211X1 ON211X1_82 ( .gnd!(gnd!), .vdd!(vdd!), .A(_840_), .B(_842_), .C(_953_), .D(_948_), .Q(_1183_) );
AN211X1 AN211X1_10 ( .gnd!(gnd!), .vdd!(vdd!), .A(_873_), .B(_875_), .C(_1183_), .D(_1182_), .Q(_1184_) );
AND5X1 AND5X1_2 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1115_), .B(_1181_), .C(_1184_), .D(_1138_), .E(_1178_), .Q(ALU_zf) );
MU2IX1 MU2IX1_104 ( .gnd!(gnd!), .vdd!(vdd!), .IN0(_1130_), .IN1(_1131_), .Q(ALU_vf), .S(_1128_) );
NA2X1 NA2X1_548 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1957_), .B(_1221__bF_buf0), .Q(_1186_) );
AND2X2 AND2X2_38 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1510_), .B(_1230__bF_buf2), .Q(_1187_) );
AND2X2 AND2X2_39 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1372_), .B(_1240__bF_buf0), .Q(_1188_) );
ON31X1 ON31X1_54 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1080_), .B(_1240__bF_buf0), .C(_1242__bF_buf3), .D(_1252__bF_buf4), .Q(_1189_) );
ON31X1 ON31X1_55 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1514_), .B(_1189_), .C(_1188_), .D(_1227__bF_buf3), .Q(_1190_) );
ON22X1 ON22X1_63 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1689_), .B(_1227__bF_buf3), .C(_1187_), .D(_1190_), .Q(_1191_) );
ON211X1 ON211X1_83 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1191_), .B(_1221__bF_buf3), .C(EXT_type_bF_buf2), .D(_1186_), .Q(_1192_) );
ON31X1 ON31X1_56 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1226__bF_buf6), .B(_1400_), .C(_1684_), .D(_1192_), .Q(_1193_) );
MU2IX1 MU2IX1_105 ( .gnd!(gnd!), .vdd!(vdd!), .IN0(_1193_), .IN1(_1161_), .Q(_1195_), .S(_952__bF_buf4) );
NA2X1 NA2X1_549 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1195_), .B(_909__bF_buf2), .Q(_1196_) );
AN211X1 AN211X1_11 ( .gnd!(gnd!), .vdd!(vdd!), .A(_984_), .B(_1327_), .C(_1160_), .D(_1330_), .Q(_1197_) );
NO2X1 NO2X1_211 ( .gnd!(gnd!), .vdd!(vdd!), .A(_995_), .B(_1526__bF_buf3), .Q(_1198_) );
ON311X1 ON311X1_7 ( .gnd!(gnd!), .vdd!(vdd!), .A(_909__bF_buf1), .B(_1197_), .C(_1198_), .D(_1143__bF_buf1), .E(_1196_), .Q(_1199_) );
NA2X1 NA2X1_550 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1163_), .B(_1112_), .Q(_1200_) );
AN211X1 AN211X1_12 ( .gnd!(gnd!), .vdd!(vdd!), .A(ALU_a_31_), .B(_1129_), .C(_1200_), .D(_1145_), .Q(_1201_) );
AN21X1 AN21X1_147 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1159_), .B(_1158_), .C(_834_), .Q(_1202_) );
ON31X1 ON31X1_57 ( .gnd!(gnd!), .vdd!(vdd!), .A(_1143__bF_buf1), .B(_1202_), .C(_1201_), .D(_1199_), .Q(ALU_r_0_) );
NO2X1 NO2X1_212 ( .gnd!(gnd!), .vdd!(vdd!), .A(CNTR_Timer_15_), .B(CNTR_Timer_14_), .Q(_2040_) );
NO2X1 NO2X1_213 ( .gnd!(gnd!), .vdd!(vdd!), .A(CNTR_Timer_8_), .B(CNTR_Timer_11_), .Q(_2041_) );
NO2X1 NO2X1_214 ( .gnd!(gnd!), .vdd!(vdd!), .A(CNTR_Timer_13_), .B(CNTR_Timer_12_), .Q(_2042_) );
NO2X1 NO2X1_215 ( .gnd!(gnd!), .vdd!(vdd!), .A(CNTR_Timer_9_), .B(CNTR_Timer_10_), .Q(_2043_) );
AND4X1 AND4X1_1 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2040_), .B(_2041_), .C(_2042_), .D(_2043_), .Q(_2044_) );
INX1 INX1_143 ( .gnd!(gnd!), .vdd!(vdd!), .A(CNTR_Timer_24_), .Q(_2045_) );
INX1 INX1_144 ( .gnd!(gnd!), .vdd!(vdd!), .A(CNTR_Timer_27_), .Q(_2046_) );
NO2X1 NO2X1_216 ( .gnd!(gnd!), .vdd!(vdd!), .A(CNTR_Timer_28_), .B(CNTR_Timer_31_), .Q(_2047_) );
NO2X1 NO2X1_217 ( .gnd!(gnd!), .vdd!(vdd!), .A(CNTR_Timer_29_), .B(CNTR_Timer_30_), .Q(_2048_) );
NO2X1 NO2X1_218 ( .gnd!(gnd!), .vdd!(vdd!), .A(CNTR_Timer_25_), .B(CNTR_Timer_26_), .Q(_2049_) );
AND5X1 AND5X1_3 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2045_), .B(_2046_), .C(_2047_), .D(_2048_), .E(_2049_), .Q(_2050_) );
NO2X1 NO2X1_219 ( .gnd!(gnd!), .vdd!(vdd!), .A(CNTR_Timer_16_), .B(CNTR_Timer_19_), .Q(_2051_) );
NO2X1 NO2X1_220 ( .gnd!(gnd!), .vdd!(vdd!), .A(CNTR_Timer_17_), .B(CNTR_Timer_18_), .Q(_2052_) );
AND2X2 AND2X2_40 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2051_), .B(_2052_), .Q(_2053_) );
NO2X1 NO2X1_221 ( .gnd!(gnd!), .vdd!(vdd!), .A(CNTR_Timer_20_), .B(CNTR_Timer_23_), .Q(_2054_) );
NO2X1 NO2X1_222 ( .gnd!(gnd!), .vdd!(vdd!), .A(CNTR_Timer_21_), .B(CNTR_Timer_22_), .Q(_2055_) );
AND2X2 AND2X2_41 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2054_), .B(_2055_), .Q(_2056_) );
AND2X2 AND2X2_42 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2053_), .B(_2056_), .Q(_2057_) );
NA3X1 NA3X1_8 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2044_), .B(_2050_), .C(_2057_), .Q(_2058_) );
NO2X1 NO2X1_223 ( .gnd!(gnd!), .vdd!(vdd!), .A(CNTR_Timer_4_), .B(CNTR_Timer_7_), .Q(_2059_) );
NO2X1 NO2X1_224 ( .gnd!(gnd!), .vdd!(vdd!), .A(CNTR_Timer_5_), .B(CNTR_Timer_6_), .Q(_2060_) );
NA2X1 NA2X1_551 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2059_), .B(_2060_), .Q(_2061_) );
NO2X1 NO2X1_225 ( .gnd!(gnd!), .vdd!(vdd!), .A(CNTR_Timer_3_), .B(CNTR_Timer_2_), .Q(_2062_) );
NA3I1X1 NA3I1X1_97 ( .gnd!(gnd!), .vdd!(vdd!), .AN(CNTR_Timer_1_), .B(CNTR_Timer_0_), .C(_2062_), .Q(_2063_) );
NO3X1 NO3X1_8 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2058_), .B(_2061_), .C(_2063_), .Q(CNTR_tif) );
MU2X1 MU2X1_202 ( .gnd!(gnd!), .vdd!(vdd!), .IN0(CNTR_gie), .IN1(_681__0_), .Q(_2039__0_), .S(CNTR_ld_uie) );
MU2X1 MU2X1_203 ( .gnd!(gnd!), .vdd!(vdd!), .IN0(CNTR_tie), .IN1(_681__1_), .Q(_2039__1_), .S(CNTR_ld_uie) );
MU2X1 MU2X1_204 ( .gnd!(gnd!), .vdd!(vdd!), .IN0(CNTR_eie), .IN1(_681__2_), .Q(_2039__2_), .S(CNTR_ld_uie) );
INX1 INX1_145 ( .gnd!(gnd!), .vdd!(vdd!), .A(_681__0_), .Q(_2064_) );
MU2IX1 MU2IX1_106 ( .gnd!(gnd!), .vdd!(vdd!), .IN0(CNTR_Cycle_0_), .IN1(_2064_), .Q(_2037__0_), .S(CNTR_ld_cycle_bF_buf5) );
NO2X1 NO2X1_226 ( .gnd!(gnd!), .vdd!(vdd!), .A(CNTR_Cycle_0_), .B(CNTR_Cycle_1_), .Q(_2065_) );
NA2X1 NA2X1_552 ( .gnd!(gnd!), .vdd!(vdd!), .A(CNTR_Cycle_0_), .B(CNTR_Cycle_1_), .Q(_2066_) );
INX1 INX1_146 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2066_), .Q(_2067_) );
NA2X1 NA2X1_553 ( .gnd!(gnd!), .vdd!(vdd!), .A(_681__1_), .B(CNTR_ld_cycle_bF_buf4), .Q(_2068_) );
ON31X1 ON31X1_58 ( .gnd!(gnd!), .vdd!(vdd!), .A(CNTR_ld_cycle_bF_buf4), .B(_2065_), .C(_2067_), .D(_2068_), .Q(_2037__1_) );
NO2X1 NO2X1_227 ( .gnd!(gnd!), .vdd!(vdd!), .A(CNTR_Cycle_2_), .B(_2067_), .Q(_2069_) );
AND2X2 AND2X2_43 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2067_), .B(CNTR_Cycle_2_), .Q(_2070_) );
NA2X1 NA2X1_554 ( .gnd!(gnd!), .vdd!(vdd!), .A(_681__2_), .B(CNTR_ld_cycle_bF_buf4), .Q(_2071_) );
ON31X1 ON31X1_59 ( .gnd!(gnd!), .vdd!(vdd!), .A(CNTR_ld_cycle_bF_buf5), .B(_2069_), .C(_2070_), .D(_2071_), .Q(_2037__2_) );
NO2X1 NO2X1_228 ( .gnd!(gnd!), .vdd!(vdd!), .A(CNTR_Cycle_3_), .B(_2070_), .Q(_2072_) );
NA2X1 NA2X1_555 ( .gnd!(gnd!), .vdd!(vdd!), .A(CNTR_Cycle_2_), .B(CNTR_Cycle_3_), .Q(_2073_) );
NO2X1 NO2X1_229 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2066_), .B(_2073_), .Q(_2074_) );
NA2X1 NA2X1_556 ( .gnd!(gnd!), .vdd!(vdd!), .A(CNTR_ld_cycle_bF_buf4), .B(_681__3_), .Q(_2075_) );
ON31X1 ON31X1_60 ( .gnd!(gnd!), .vdd!(vdd!), .A(CNTR_ld_cycle_bF_buf4), .B(_2074_), .C(_2072_), .D(_2075_), .Q(_2037__3_) );
INX1 INX1_147 ( .gnd!(gnd!), .vdd!(vdd!), .A(CNTR_ld_cycle_bF_buf5), .Q(_2076_) );
INX1 INX1_148 ( .gnd!(gnd!), .vdd!(vdd!), .A(_681__4_), .Q(_2077_) );
NO2X1 NO2X1_230 ( .gnd!(gnd!), .vdd!(vdd!), .A(CNTR_Cycle_4_), .B(_2074_), .Q(_2078_) );
NA2X1 NA2X1_557 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2074_), .B(CNTR_Cycle_4_), .Q(_2079_) );
NA2X1 NA2X1_558 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2079_), .B(_2076_), .Q(_2080_) );
ON22X1 ON22X1_64 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2080_), .B(_2078_), .C(_2076_), .D(_2077_), .Q(_2037__4_) );
INX1 INX1_149 ( .gnd!(gnd!), .vdd!(vdd!), .A(CNTR_Cycle_5_), .Q(_2081_) );
NO2X1 NO2X1_231 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2081_), .B(_2079_), .Q(_2082_) );
AND2X2 AND2X2_44 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2079_), .B(_2081_), .Q(_2083_) );
NA2X1 NA2X1_559 ( .gnd!(gnd!), .vdd!(vdd!), .A(CNTR_ld_cycle_bF_buf5), .B(_681__5_), .Q(_2084_) );
ON31X1 ON31X1_61 ( .gnd!(gnd!), .vdd!(vdd!), .A(CNTR_ld_cycle_bF_buf5), .B(_2082_), .C(_2083_), .D(_2084_), .Q(_2037__5_) );
NO2X1 NO2X1_232 ( .gnd!(gnd!), .vdd!(vdd!), .A(CNTR_Cycle_6_), .B(_2082_), .Q(_2085_) );
AND2X2 AND2X2_45 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2082_), .B(CNTR_Cycle_6_), .Q(_2086_) );
NA2X1 NA2X1_560 ( .gnd!(gnd!), .vdd!(vdd!), .A(CNTR_ld_cycle_bF_buf5), .B(_681__6_), .Q(_2087_) );
ON31X1 ON31X1_62 ( .gnd!(gnd!), .vdd!(vdd!), .A(CNTR_ld_cycle_bF_buf5), .B(_2085_), .C(_2086_), .D(_2087_), .Q(_2037__6_) );
INX1 INX1_150 ( .gnd!(gnd!), .vdd!(vdd!), .A(_681__7_), .Q(_2088_) );
NO2X1 NO2X1_233 ( .gnd!(gnd!), .vdd!(vdd!), .A(CNTR_Cycle_7_), .B(_2086_), .Q(_2089_) );
AND4X1 AND4X1_2 ( .gnd!(gnd!), .vdd!(vdd!), .A(CNTR_Cycle_4_), .B(CNTR_Cycle_5_), .C(CNTR_Cycle_6_), .D(CNTR_Cycle_7_), .Q(_2090_) );
NA2X1 NA2X1_561 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2074_), .B(_2090_), .Q(_2091_) );
NA2X1 NA2X1_562 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2091_), .B(_2076_), .Q(_2092_) );
ON22X1 ON22X1_65 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2089_), .B(_2092_), .C(_2076_), .D(_2088_), .Q(_2037__7_) );
NO2I1X1 NO2I1X1_37 ( .gnd!(gnd!), .vdd!(vdd!), .AN(CNTR_Cycle_8_), .B(_2091_), .Q(_2093_) );
AND2X2 AND2X2_46 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2074_), .B(_2090_), .Q(_2094_) );
NO2X1 NO2X1_234 ( .gnd!(gnd!), .vdd!(vdd!), .A(CNTR_Cycle_8_), .B(_2094_), .Q(_2095_) );
NA2X1 NA2X1_563 ( .gnd!(gnd!), .vdd!(vdd!), .A(CNTR_ld_cycle_bF_buf6), .B(_681__8_), .Q(_2096_) );
ON31X1 ON31X1_63 ( .gnd!(gnd!), .vdd!(vdd!), .A(CNTR_ld_cycle_bF_buf6), .B(_2093_), .C(_2095_), .D(_2096_), .Q(_2037__8_) );
INX1 INX1_151 ( .gnd!(gnd!), .vdd!(vdd!), .A(_681__9_), .Q(_2097_) );
NO2X1 NO2X1_235 ( .gnd!(gnd!), .vdd!(vdd!), .A(CNTR_Cycle_9_), .B(_2093_), .Q(_2098_) );
NA2X1 NA2X1_564 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2093_), .B(CNTR_Cycle_9_), .Q(_2099_) );
NA2X1 NA2X1_565 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2099_), .B(_2076_), .Q(_2100_) );
ON22X1 ON22X1_66 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2100_), .B(_2098_), .C(_2076_), .D(_2097_), .Q(_2037__9_) );
INX1 INX1_152 ( .gnd!(gnd!), .vdd!(vdd!), .A(CNTR_Cycle_10_), .Q(_2101_) );
NO2X1 NO2X1_236 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2101_), .B(_2099_), .Q(_2102_) );
AND2X2 AND2X2_47 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2099_), .B(_2101_), .Q(_2103_) );
NA2X1 NA2X1_566 ( .gnd!(gnd!), .vdd!(vdd!), .A(CNTR_ld_cycle_bF_buf6), .B(_681__10_), .Q(_2104_) );
ON31X1 ON31X1_64 ( .gnd!(gnd!), .vdd!(vdd!), .A(CNTR_ld_cycle_bF_buf6), .B(_2102_), .C(_2103_), .D(_2104_), .Q(_2037__10_) );
NA2X1 NA2X1_567 ( .gnd!(gnd!), .vdd!(vdd!), .A(CNTR_ld_cycle_bF_buf3), .B(_681__11_), .Q(_2105_) );
NO2X1 NO2X1_237 ( .gnd!(gnd!), .vdd!(vdd!), .A(CNTR_Cycle_11_), .B(_2102_), .Q(_2106_) );
AND4X1 AND4X1_3 ( .gnd!(gnd!), .vdd!(vdd!), .A(CNTR_Cycle_8_), .B(CNTR_Cycle_9_), .C(CNTR_Cycle_10_), .D(CNTR_Cycle_11_), .Q(_2107_) );
NA2X1 NA2X1_568 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2094_), .B(_2107_), .Q(_2108_) );
NA2X1 NA2X1_569 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2108_), .B(_2076_), .Q(_2109_) );
ON21X1 ON21X1_281 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2106_), .B(_2109_), .C(_2105_), .Q(_2037__11_) );
INX1 INX1_153 ( .gnd!(gnd!), .vdd!(vdd!), .A(CNTR_Cycle_12_), .Q(_2110_) );
NO2X1 NO2X1_238 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2110_), .B(_2108_), .Q(_2111_) );
AND2X2 AND2X2_48 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2108_), .B(_2110_), .Q(_2112_) );
NA2X1 NA2X1_570 ( .gnd!(gnd!), .vdd!(vdd!), .A(CNTR_ld_cycle_bF_buf3), .B(_681__12_), .Q(_2113_) );
ON31X1 ON31X1_65 ( .gnd!(gnd!), .vdd!(vdd!), .A(CNTR_ld_cycle_bF_buf3), .B(_2111_), .C(_2112_), .D(_2113_), .Q(_2037__12_) );
NA2X1 NA2X1_571 ( .gnd!(gnd!), .vdd!(vdd!), .A(CNTR_ld_cycle_bF_buf3), .B(_681__13_), .Q(_2114_) );
NO2X1 NO2X1_239 ( .gnd!(gnd!), .vdd!(vdd!), .A(CNTR_Cycle_13_), .B(_2111_), .Q(_2115_) );
AND4X1 AND4X1_4 ( .gnd!(gnd!), .vdd!(vdd!), .A(CNTR_Cycle_12_), .B(CNTR_Cycle_13_), .C(_2107_), .D(_2094_), .Q(_2116_) );
ON31X1 ON31X1_66 ( .gnd!(gnd!), .vdd!(vdd!), .A(CNTR_ld_cycle_bF_buf3), .B(_2116_), .C(_2115_), .D(_2114_), .Q(_2037__13_) );
NA2X1 NA2X1_572 ( .gnd!(gnd!), .vdd!(vdd!), .A(CNTR_ld_cycle_bF_buf3), .B(_681__14_), .Q(_2117_) );
NO2X1 NO2X1_240 ( .gnd!(gnd!), .vdd!(vdd!), .A(CNTR_Cycle_14_), .B(_2116_), .Q(_2118_) );
AND2X2 AND2X2_49 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2116_), .B(CNTR_Cycle_14_), .Q(_2119_) );
ON31X1 ON31X1_67 ( .gnd!(gnd!), .vdd!(vdd!), .A(CNTR_ld_cycle_bF_buf3), .B(_2118_), .C(_2119_), .D(_2117_), .Q(_2037__14_) );
NA2X1 NA2X1_573 ( .gnd!(gnd!), .vdd!(vdd!), .A(CNTR_Cycle_12_), .B(CNTR_Cycle_13_), .Q(_2120_) );
NO2X1 NO2X1_241 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2120_), .B(_2108_), .Q(_2121_) );
NA2X1 NA2X1_574 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2121_), .B(CNTR_Cycle_14_), .Q(_2122_) );
NA2X1 NA2X1_575 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2122_), .B(CNTR_Cycle_15_), .Q(_2123_) );
NA3I1X1 NA3I1X1_98 ( .gnd!(gnd!), .vdd!(vdd!), .AN(CNTR_Cycle_15_), .B(CNTR_Cycle_14_), .C(_2121_), .Q(_2124_) );
NO2X1 NO2X1_242 ( .gnd!(gnd!), .vdd!(vdd!), .A(_681__15_), .B(_2076_), .Q(_2125_) );
AN31X1 AN31X1_62 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2076_), .B(_2124_), .C(_2123_), .D(_2125_), .Q(_2037__15_) );
INX1 INX1_154 ( .gnd!(gnd!), .vdd!(vdd!), .A(_681__16_), .Q(_2126_) );
AND2X2 AND2X2_50 ( .gnd!(gnd!), .vdd!(vdd!), .A(CNTR_Cycle_14_), .B(CNTR_Cycle_15_), .Q(_2127_) );
NA3I1X1 NA3I1X1_99 ( .gnd!(gnd!), .vdd!(vdd!), .AN(_2120_), .B(_2127_), .C(_2107_), .Q(_2128_) );
NO2X1 NO2X1_243 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2091_), .B(_2128_), .Q(_2129_) );
EN2X1 EN2X1_11 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2129_), .B(CNTR_Cycle_16_), .Q(_2130_) );
MU2IX1 MU2IX1_107 ( .gnd!(gnd!), .vdd!(vdd!), .IN0(_2130_), .IN1(_2126_), .Q(_2037__16_), .S(CNTR_ld_cycle_bF_buf2) );
NA2X1 NA2X1_576 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2129_), .B(CNTR_Cycle_16_), .Q(_2131_) );
NA2I1X1 NA2I1X1_74 ( .gnd!(gnd!), .vdd!(vdd!), .AN(CNTR_Cycle_17_), .B(_2131_), .Q(_2132_) );
AND2X2 AND2X2_51 ( .gnd!(gnd!), .vdd!(vdd!), .A(CNTR_Cycle_16_), .B(CNTR_Cycle_17_), .Q(_2133_) );
NA2X1 NA2X1_577 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2129_), .B(_2133_), .Q(_2134_) );
AND2X2 AND2X2_52 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2134_), .B(_2076_), .Q(_2135_) );
AO22X2 AO22X2_29 ( .gnd!(gnd!), .vdd!(vdd!), .A(CNTR_ld_cycle_bF_buf6), .B(_681__17_), .C(_2135_), .D(_2132_), .Q(_2037__17_) );
INX1 INX1_155 ( .gnd!(gnd!), .vdd!(vdd!), .A(CNTR_Cycle_18_), .Q(_2136_) );
NO2X1 NO2X1_244 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2136_), .B(_2134_), .Q(_2137_) );
AND2X2 AND2X2_53 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2134_), .B(_2136_), .Q(_2138_) );
NA2X1 NA2X1_578 ( .gnd!(gnd!), .vdd!(vdd!), .A(CNTR_ld_cycle_bF_buf0), .B(_681__18_), .Q(_2139_) );
ON31X1 ON31X1_68 ( .gnd!(gnd!), .vdd!(vdd!), .A(CNTR_ld_cycle_bF_buf0), .B(_2137_), .C(_2138_), .D(_2139_), .Q(_2037__18_) );
NA2X1 NA2X1_579 ( .gnd!(gnd!), .vdd!(vdd!), .A(CNTR_ld_cycle_bF_buf2), .B(_681__19_), .Q(_2140_) );
NO2X1 NO2X1_245 ( .gnd!(gnd!), .vdd!(vdd!), .A(CNTR_Cycle_19_), .B(_2137_), .Q(_2141_) );
AND3X4 AND3X4_8 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2133_), .B(CNTR_Cycle_18_), .C(CNTR_Cycle_19_), .Q(_2142_) );
AND2X2 AND2X2_54 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2129_), .B(_2142_), .Q(_2143_) );
ON31X1 ON31X1_69 ( .gnd!(gnd!), .vdd!(vdd!), .A(CNTR_ld_cycle_bF_buf2), .B(_2143_), .C(_2141_), .D(_2140_), .Q(_2037__19_) );
AND2X2 AND2X2_55 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2143_), .B(CNTR_Cycle_20_), .Q(_2144_) );
NO2X1 NO2X1_246 ( .gnd!(gnd!), .vdd!(vdd!), .A(CNTR_Cycle_20_), .B(_2143_), .Q(_2145_) );
NA2X1 NA2X1_580 ( .gnd!(gnd!), .vdd!(vdd!), .A(CNTR_ld_cycle_bF_buf2), .B(_681__20_), .Q(_2146_) );
ON31X1 ON31X1_70 ( .gnd!(gnd!), .vdd!(vdd!), .A(CNTR_ld_cycle_bF_buf2), .B(_2145_), .C(_2144_), .D(_2146_), .Q(_2037__20_) );
NA2X1 NA2X1_581 ( .gnd!(gnd!), .vdd!(vdd!), .A(CNTR_ld_cycle_bF_buf2), .B(_681__21_), .Q(_2147_) );
AN31X1 AN31X1_63 ( .gnd!(gnd!), .vdd!(vdd!), .A(CNTR_Cycle_20_), .B(_2142_), .C(_2129_), .D(CNTR_Cycle_21_), .Q(_2148_) );
AND4X1 AND4X1_5 ( .gnd!(gnd!), .vdd!(vdd!), .A(CNTR_Cycle_20_), .B(CNTR_Cycle_21_), .C(_2142_), .D(_2129_), .Q(_2149_) );
ON31X1 ON31X1_71 ( .gnd!(gnd!), .vdd!(vdd!), .A(CNTR_ld_cycle_bF_buf2), .B(_2148_), .C(_2149_), .D(_2147_), .Q(_2037__21_) );
NA2X1 NA2X1_582 ( .gnd!(gnd!), .vdd!(vdd!), .A(CNTR_ld_cycle_bF_buf6), .B(_681__22_), .Q(_2150_) );
NO2X1 NO2X1_247 ( .gnd!(gnd!), .vdd!(vdd!), .A(CNTR_Cycle_22_), .B(_2149_), .Q(_2151_) );
AND5X1 AND5X1_4 ( .gnd!(gnd!), .vdd!(vdd!), .A(CNTR_Cycle_20_), .B(CNTR_Cycle_21_), .C(CNTR_Cycle_22_), .D(_2142_), .E(_2129_), .Q(_2152_) );
ON31X1 ON31X1_72 ( .gnd!(gnd!), .vdd!(vdd!), .A(CNTR_ld_cycle_bF_buf6), .B(_2152_), .C(_2151_), .D(_2150_), .Q(_2037__22_) );
NA2X1 NA2X1_583 ( .gnd!(gnd!), .vdd!(vdd!), .A(CNTR_ld_cycle_bF_buf0), .B(_681__23_), .Q(_2153_) );
NO2X1 NO2X1_248 ( .gnd!(gnd!), .vdd!(vdd!), .A(CNTR_Cycle_23_), .B(_2152_), .Q(_2154_) );
AND4X1 AND4X1_6 ( .gnd!(gnd!), .vdd!(vdd!), .A(CNTR_Cycle_20_), .B(CNTR_Cycle_21_), .C(CNTR_Cycle_22_), .D(CNTR_Cycle_23_), .Q(_2155_) );
AND4X1 AND4X1_7 ( .gnd!(gnd!), .vdd!(vdd!), .A(CNTR_Cycle_18_), .B(CNTR_Cycle_19_), .C(_2133_), .D(_2155_), .Q(_2156_) );
AND2X2 AND2X2_56 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2129_), .B(_2156_), .Q(_2157_) );
ON31X1 ON31X1_73 ( .gnd!(gnd!), .vdd!(vdd!), .A(CNTR_ld_cycle_bF_buf0), .B(_2157_), .C(_2154_), .D(_2153_), .Q(_2037__23_) );
AND2X2 AND2X2_57 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2157_), .B(CNTR_Cycle_24_), .Q(_2158_) );
NO2X1 NO2X1_249 ( .gnd!(gnd!), .vdd!(vdd!), .A(CNTR_Cycle_24_), .B(_2157_), .Q(_2159_) );
NA2X1 NA2X1_584 ( .gnd!(gnd!), .vdd!(vdd!), .A(CNTR_ld_cycle_bF_buf0), .B(_681__24_), .Q(_2160_) );
ON31X1 ON31X1_74 ( .gnd!(gnd!), .vdd!(vdd!), .A(CNTR_ld_cycle_bF_buf0), .B(_2159_), .C(_2158_), .D(_2160_), .Q(_2037__24_) );
NA2X1 NA2X1_585 ( .gnd!(gnd!), .vdd!(vdd!), .A(CNTR_ld_cycle_bF_buf1), .B(_681__25_), .Q(_2161_) );
AN31X1 AN31X1_64 ( .gnd!(gnd!), .vdd!(vdd!), .A(CNTR_Cycle_24_), .B(_2156_), .C(_2129_), .D(CNTR_Cycle_25_), .Q(_2162_) );
AND2X2 AND2X2_58 ( .gnd!(gnd!), .vdd!(vdd!), .A(CNTR_Cycle_24_), .B(CNTR_Cycle_25_), .Q(_2163_) );
AND2X2 AND2X2_59 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2157_), .B(_2163_), .Q(_2164_) );
ON31X1 ON31X1_75 ( .gnd!(gnd!), .vdd!(vdd!), .A(CNTR_ld_cycle_bF_buf0), .B(_2162_), .C(_2164_), .D(_2161_), .Q(_2037__25_) );
INX1 INX1_156 ( .gnd!(gnd!), .vdd!(vdd!), .A(_681__26_), .Q(_2165_) );
AN31X1 AN31X1_65 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2156_), .B(_2163_), .C(_2129_), .D(CNTR_Cycle_26_), .Q(_2166_) );
AND2X2 AND2X2_60 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2163_), .B(CNTR_Cycle_26_), .Q(_2167_) );
NA2X1 NA2X1_586 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2157_), .B(_2167_), .Q(_2168_) );
NA2X1 NA2X1_587 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2168_), .B(_2076_), .Q(_2169_) );
ON22X1 ON22X1_67 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2169_), .B(_2166_), .C(_2076_), .D(_2165_), .Q(_2037__26_) );
AN31X1 AN31X1_66 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2156_), .B(_2167_), .C(_2129_), .D(CNTR_Cycle_27_), .Q(_2170_) );
AND4X1 AND4X1_8 ( .gnd!(gnd!), .vdd!(vdd!), .A(CNTR_Cycle_27_), .B(_2156_), .C(_2167_), .D(_2129_), .Q(_2171_) );
NA2X1 NA2X1_588 ( .gnd!(gnd!), .vdd!(vdd!), .A(CNTR_ld_cycle_bF_buf4), .B(_681__27_), .Q(_2172_) );
ON31X1 ON31X1_76 ( .gnd!(gnd!), .vdd!(vdd!), .A(CNTR_ld_cycle_bF_buf1), .B(_2170_), .C(_2171_), .D(_2172_), .Q(_2037__27_) );
NO2X1 NO2X1_250 ( .gnd!(gnd!), .vdd!(vdd!), .A(CNTR_Cycle_28_), .B(_2171_), .Q(_2173_) );
AND3X4 AND3X4_9 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2163_), .B(CNTR_Cycle_26_), .C(CNTR_Cycle_27_), .Q(_2174_) );
NA3X1 NA3X1_9 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2156_), .B(_2174_), .C(_2129_), .Q(_2175_) );
NO2I1X1 NO2I1X1_38 ( .gnd!(gnd!), .vdd!(vdd!), .AN(CNTR_Cycle_28_), .B(_2175_), .Q(_2176_) );
NA2X1 NA2X1_589 ( .gnd!(gnd!), .vdd!(vdd!), .A(CNTR_ld_cycle_bF_buf1), .B(_681__28_), .Q(_2177_) );
ON31X1 ON31X1_77 ( .gnd!(gnd!), .vdd!(vdd!), .A(CNTR_ld_cycle_bF_buf1), .B(_2176_), .C(_2173_), .D(_2177_), .Q(_2037__28_) );
NO2X1 NO2X1_251 ( .gnd!(gnd!), .vdd!(vdd!), .A(CNTR_Cycle_29_), .B(_2176_), .Q(_2178_) );
AND2X2 AND2X2_61 ( .gnd!(gnd!), .vdd!(vdd!), .A(CNTR_Cycle_28_), .B(CNTR_Cycle_29_), .Q(_2179_) );
NO2I1X1 NO2I1X1_39 ( .gnd!(gnd!), .vdd!(vdd!), .AN(_2179_), .B(_2175_), .Q(_2180_) );
NA2X1 NA2X1_590 ( .gnd!(gnd!), .vdd!(vdd!), .A(CNTR_ld_cycle_bF_buf1), .B(_681__29_), .Q(_2181_) );
ON31X1 ON31X1_78 ( .gnd!(gnd!), .vdd!(vdd!), .A(CNTR_ld_cycle_bF_buf1), .B(_2180_), .C(_2178_), .D(_2181_), .Q(_2037__29_) );
NO2X1 NO2X1_252 ( .gnd!(gnd!), .vdd!(vdd!), .A(CNTR_Cycle_30_), .B(_2180_), .Q(_2182_) );
AND5X1 AND5X1_5 ( .gnd!(gnd!), .vdd!(vdd!), .A(CNTR_Cycle_30_), .B(_2174_), .C(_2179_), .D(_2156_), .E(_2129_), .Q(_2183_) );
NA2X1 NA2X1_591 ( .gnd!(gnd!), .vdd!(vdd!), .A(CNTR_ld_cycle_bF_buf4), .B(_681__30_), .Q(_2184_) );
ON31X1 ON31X1_79 ( .gnd!(gnd!), .vdd!(vdd!), .A(CNTR_ld_cycle_bF_buf1), .B(_2183_), .C(_2182_), .D(_2184_), .Q(_2037__30_) );
INX1 INX1_157 ( .gnd!(gnd!), .vdd!(vdd!), .A(_681__31_), .Q(_2185_) );
AND2X2 AND2X2_62 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2183_), .B(CNTR_Cycle_31_), .Q(_2186_) );
ON21X1 ON21X1_282 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2183_), .B(CNTR_Cycle_31_), .C(_2076_), .Q(_2187_) );
ON22X1 ON22X1_68 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2186_), .B(_2187_), .C(_2076_), .D(_2185_), .Q(_2037__31_) );
INX1 INX1_158 ( .gnd!(gnd!), .vdd!(vdd!), .A(CNTR_ld_timer_bF_buf2), .Q(_2188_) );
NO2X1 NO2X1_253 ( .gnd!(gnd!), .vdd!(vdd!), .A(CNTR_Timer_0_), .B(CNTR_Timer_1_), .Q(_2189_) );
NA2X1 NA2X1_592 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2062_), .B(_2189_), .Q(_2190_) );
OR2X2 OR2X2_13 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2061_), .B(_2190_), .Q(_2191_) );
ON21X1 ON21X1_283 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2058_), .B(_2191_), .C(_2188_), .Q(_2192_) );
ON22X1 ON22X1_69 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2192_), .B(CNTR_Timer_0_), .C(_2064_), .D(_2188_), .Q(_2038__0_) );
NO2X1 NO2X1_254 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2061_), .B(_2190_), .Q(_2193_) );
AND2X2 AND2X2_63 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2193_), .B(_2044_), .Q(_2194_) );
AN31X1 AN31X1_67 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2050_), .B(_2057_), .C(_2194_), .D(CNTR_ld_timer_bF_buf0), .Q(_2195_) );
EN2X1 EN2X1_12 ( .gnd!(gnd!), .vdd!(vdd!), .A(CNTR_Timer_0_), .B(CNTR_Timer_1_), .Q(_2196_) );
AO22X2 AO22X2_30 ( .gnd!(gnd!), .vdd!(vdd!), .A(_681__1_), .B(CNTR_ld_timer_bF_buf4), .C(_2195__bF_buf3), .D(_2196_), .Q(_2038__1_) );
NA2I1X1 NA2I1X1_75 ( .gnd!(gnd!), .vdd!(vdd!), .AN(CNTR_Timer_2_), .B(_2189_), .Q(_2197_) );
NA2I1X1 NA2I1X1_76 ( .gnd!(gnd!), .vdd!(vdd!), .AN(_2189_), .B(CNTR_Timer_2_), .Q(_2198_) );
NA2X1 NA2X1_593 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2198_), .B(_2197_), .Q(_2199_) );
AO22X2 AO22X2_31 ( .gnd!(gnd!), .vdd!(vdd!), .A(_681__2_), .B(CNTR_ld_timer_bF_buf4), .C(_2195__bF_buf3), .D(_2199_), .Q(_2038__2_) );
NA2X1 NA2X1_594 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2197_), .B(CNTR_Timer_3_), .Q(_2200_) );
NA2X1 NA2X1_595 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2200_), .B(_2190_), .Q(_2201_) );
AO22X2 AO22X2_32 ( .gnd!(gnd!), .vdd!(vdd!), .A(_681__3_), .B(CNTR_ld_timer_bF_buf4), .C(_2195__bF_buf3), .D(_2201_), .Q(_2038__3_) );
INX1 INX1_159 ( .gnd!(gnd!), .vdd!(vdd!), .A(CNTR_Timer_4_), .Q(_2202_) );
EN2X1 EN2X1_13 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2190_), .B(_2202_), .Q(_2203_) );
ON22X1 ON22X1_70 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2192_), .B(_2203_), .C(_2077_), .D(_2188_), .Q(_2038__4_) );
NA2I1X1 NA2I1X1_77 ( .gnd!(gnd!), .vdd!(vdd!), .AN(_2190_), .B(_2202_), .Q(_2204_) );
NA2X1 NA2X1_596 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2204_), .B(CNTR_Timer_5_), .Q(_2205_) );
OR2X2 OR2X2_14 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2204_), .B(CNTR_Timer_5_), .Q(_2206_) );
NA2X1 NA2X1_597 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2206_), .B(_2205_), .Q(_2207_) );
AO22X2 AO22X2_33 ( .gnd!(gnd!), .vdd!(vdd!), .A(_681__5_), .B(CNTR_ld_timer_bF_buf4), .C(_2195__bF_buf3), .D(_2207_), .Q(_2038__5_) );
NA2X1 NA2X1_598 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2206_), .B(CNTR_Timer_6_), .Q(_2208_) );
NA2I1X1 NA2I1X1_78 ( .gnd!(gnd!), .vdd!(vdd!), .AN(_2204_), .B(_2060_), .Q(_2209_) );
NA2X1 NA2X1_599 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2208_), .B(_2209_), .Q(_2210_) );
AO22X2 AO22X2_34 ( .gnd!(gnd!), .vdd!(vdd!), .A(_681__6_), .B(CNTR_ld_timer_bF_buf4), .C(_2210_), .D(_2195__bF_buf3), .Q(_2038__6_) );
AN21X1 AN21X1_148 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2209_), .B(CNTR_Timer_7_), .C(_2193_), .Q(_2211_) );
ON22X1 ON22X1_71 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2192_), .B(_2211_), .C(_2088_), .D(_2188_), .Q(_2038__7_) );
NA2X1 NA2X1_600 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2191_), .B(CNTR_Timer_8_), .Q(_2212_) );
INX1 INX1_160 ( .gnd!(gnd!), .vdd!(vdd!), .A(CNTR_Timer_8_), .Q(_2213_) );
NA2X1 NA2X1_601 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2193_), .B(_2213_), .Q(_2214_) );
NA2X1 NA2X1_602 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2212_), .B(_2214_), .Q(_2215_) );
AO22X2 AO22X2_35 ( .gnd!(gnd!), .vdd!(vdd!), .A(_681__8_), .B(CNTR_ld_timer_bF_buf4), .C(_2195__bF_buf3), .D(_2215_), .Q(_2038__8_) );
NO2X1 NO2X1_255 ( .gnd!(gnd!), .vdd!(vdd!), .A(CNTR_Timer_8_), .B(_2191_), .Q(_2216_) );
EN2X1 EN2X1_14 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2216_), .B(CNTR_Timer_9_), .Q(_2217_) );
ON22X1 ON22X1_72 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2217_), .B(_2192_), .C(_2097_), .D(_2188_), .Q(_2038__9_) );
INX1 INX1_161 ( .gnd!(gnd!), .vdd!(vdd!), .A(CNTR_Timer_10_), .Q(_2218_) );
NO2X1 NO2X1_256 ( .gnd!(gnd!), .vdd!(vdd!), .A(CNTR_Timer_9_), .B(_2214_), .Q(_2219_) );
EO2X1 EO2X1_1 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2218_), .B(_2219_), .Q(_2220_) );
NA2X1 NA2X1_603 ( .gnd!(gnd!), .vdd!(vdd!), .A(_681__10_), .B(CNTR_ld_timer_bF_buf2), .Q(_2221_) );
ON21X1 ON21X1_284 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2220_), .B(_2192_), .C(_2221_), .Q(_2038__10_) );
INX1 INX1_162 ( .gnd!(gnd!), .vdd!(vdd!), .A(CNTR_Timer_11_), .Q(_2222_) );
AN31X1 AN31X1_68 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2213_), .B(_2043_), .C(_2193_), .D(_2222_), .Q(_2223_) );
AND3X4 AND3X4_10 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2216_), .B(_2222_), .C(_2043_), .Q(_2224_) );
NO2X1 NO2X1_257 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2223_), .B(_2224_), .Q(_2225_) );
NA2X1 NA2X1_604 ( .gnd!(gnd!), .vdd!(vdd!), .A(_681__11_), .B(CNTR_ld_timer_bF_buf2), .Q(_2226_) );
ON21X1 ON21X1_285 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2225_), .B(_2192_), .C(_2226_), .Q(_2038__11_) );
NO2X1 NO2X1_258 ( .gnd!(gnd!), .vdd!(vdd!), .A(CNTR_Timer_11_), .B(CNTR_Timer_12_), .Q(_2227_) );
AND4X1 AND4X1_9 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2213_), .B(_2227_), .C(_2043_), .D(_2193_), .Q(_2228_) );
INX1 INX1_163 ( .gnd!(gnd!), .vdd!(vdd!), .A(CNTR_Timer_12_), .Q(_2229_) );
AN31X1 AN31X1_69 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2222_), .B(_2043_), .C(_2216_), .D(_2229_), .Q(_2230_) );
ON21X1 ON21X1_286 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2230_), .B(_2228_), .C(_2195__bF_buf0), .Q(_2231_) );
NA2X1 NA2X1_605 ( .gnd!(gnd!), .vdd!(vdd!), .A(_681__12_), .B(CNTR_ld_timer_bF_buf0), .Q(_2232_) );
NA2X1 NA2X1_606 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2231_), .B(_2232_), .Q(_2038__12_) );
INX1 INX1_164 ( .gnd!(gnd!), .vdd!(vdd!), .A(CNTR_Timer_13_), .Q(_2233_) );
NO2X1 NO2X1_259 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2233_), .B(_2228_), .Q(_2234_) );
AND2X2 AND2X2_64 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2228_), .B(_2233_), .Q(_2235_) );
ON21X1 ON21X1_287 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2235_), .B(_2234_), .C(_2195__bF_buf1), .Q(_2236_) );
NA2X1 NA2X1_607 ( .gnd!(gnd!), .vdd!(vdd!), .A(_681__13_), .B(CNTR_ld_timer_bF_buf0), .Q(_2237_) );
NA2X1 NA2X1_608 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2236_), .B(_2237_), .Q(_2038__13_) );
INX1 INX1_165 ( .gnd!(gnd!), .vdd!(vdd!), .A(CNTR_Timer_14_), .Q(_2238_) );
AN21X1 AN21X1_149 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2228_), .B(_2233_), .C(_2238_), .Q(_2239_) );
NO2X1 NO2X1_260 ( .gnd!(gnd!), .vdd!(vdd!), .A(CNTR_Timer_13_), .B(CNTR_Timer_14_), .Q(_2240_) );
AND5X1 AND5X1_6 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2213_), .B(_2227_), .C(_2240_), .D(_2043_), .E(_2193_), .Q(_2241_) );
ON21X1 ON21X1_288 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2239_), .B(_2241_), .C(_2195__bF_buf0), .Q(_2242_) );
NA2X1 NA2X1_609 ( .gnd!(gnd!), .vdd!(vdd!), .A(_681__14_), .B(CNTR_ld_timer_bF_buf2), .Q(_2244_) );
NA2X1 NA2X1_610 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2242_), .B(_2244_), .Q(_2038__14_) );
INX1 INX1_166 ( .gnd!(gnd!), .vdd!(vdd!), .A(CNTR_Timer_15_), .Q(_2245_) );
NA2X1 NA2X1_611 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2193_), .B(_2044_), .Q(_2246_) );
ON21X1 ON21X1_289 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2241_), .B(_2245_), .C(_2246_), .Q(_2247_) );
AO22X2 AO22X2_36 ( .gnd!(gnd!), .vdd!(vdd!), .A(_681__15_), .B(CNTR_ld_timer_bF_buf0), .C(_2195__bF_buf0), .D(_2247_), .Q(_2038__15_) );
NA3I1X1 NA3I1X1_100 ( .gnd!(gnd!), .vdd!(vdd!), .AN(CNTR_Timer_16_), .B(_2044_), .C(_2193_), .Q(_2248_) );
NA2X1 NA2X1_612 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2246_), .B(CNTR_Timer_16_), .Q(_2249_) );
AND2X2 AND2X2_65 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2249_), .B(_2248_), .Q(_2250_) );
ON22X1 ON22X1_73 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2192_), .B(_2250_), .C(_2126_), .D(_2188_), .Q(_2038__16_) );
AND2X2 AND2X2_66 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2248_), .B(CNTR_Timer_17_), .Q(_2251_) );
NO2X1 NO2X1_261 ( .gnd!(gnd!), .vdd!(vdd!), .A(CNTR_Timer_17_), .B(_2248_), .Q(_2252_) );
ON21X1 ON21X1_290 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2251_), .B(_2252_), .C(_2195__bF_buf2), .Q(_2253_) );
NA2X1 NA2X1_613 ( .gnd!(gnd!), .vdd!(vdd!), .A(_681__17_), .B(CNTR_ld_timer_bF_buf3), .Q(_2254_) );
NA2X1 NA2X1_614 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2253_), .B(_2254_), .Q(_2038__17_) );
ON21X1 ON21X1_291 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2248_), .B(CNTR_Timer_17_), .C(CNTR_Timer_18_), .Q(_2255_) );
NA2I1X1 NA2I1X1_79 ( .gnd!(gnd!), .vdd!(vdd!), .AN(_2248_), .B(_2052_), .Q(_2256_) );
NA2X1 NA2X1_615 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2256_), .B(_2255_), .Q(_2257_) );
AO22X2 AO22X2_37 ( .gnd!(gnd!), .vdd!(vdd!), .A(_681__18_), .B(CNTR_ld_timer_bF_buf3), .C(_2257_), .D(_2195__bF_buf2), .Q(_2038__18_) );
ON31X1 ON31X1_80 ( .gnd!(gnd!), .vdd!(vdd!), .A(CNTR_Timer_17_), .B(CNTR_Timer_18_), .C(_2248_), .D(CNTR_Timer_19_), .Q(_2258_) );
OR2X2 OR2X2_15 ( .gnd!(gnd!), .vdd!(vdd!), .A(CNTR_Timer_8_), .B(CNTR_Timer_11_), .Q(_2259_) );
NA3X1 NA3X1_10 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2040_), .B(_2042_), .C(_2043_), .Q(_2260_) );
NA2X1 NA2X1_616 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2051_), .B(_2052_), .Q(_2261_) );
NO3X1 NO3X1_9 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2260_), .B(_2261_), .C(_2259_), .Q(_2262_) );
NA2X1 NA2X1_617 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2262_), .B(_2193_), .Q(_2263_) );
NA2X1 NA2X1_618 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2258_), .B(_2263_), .Q(_2264_) );
AO22X2 AO22X2_38 ( .gnd!(gnd!), .vdd!(vdd!), .A(_681__19_), .B(CNTR_ld_timer_bF_buf3), .C(_2264_), .D(_2195__bF_buf2), .Q(_2038__19_) );
NO2X1 NO2X1_262 ( .gnd!(gnd!), .vdd!(vdd!), .A(CNTR_Timer_20_), .B(_2263_), .Q(_2265_) );
INX1 INX1_167 ( .gnd!(gnd!), .vdd!(vdd!), .A(CNTR_Timer_20_), .Q(_2266_) );
NO2X1 NO2X1_263 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2261_), .B(_2246_), .Q(_2267_) );
NO2X1 NO2X1_264 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2266_), .B(_2267_), .Q(_2268_) );
ON21X1 ON21X1_292 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2268_), .B(_2265_), .C(_2195__bF_buf2), .Q(_2269_) );
NA2X1 NA2X1_619 ( .gnd!(gnd!), .vdd!(vdd!), .A(_681__20_), .B(CNTR_ld_timer_bF_buf3), .Q(_2270_) );
NA2X1 NA2X1_620 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2269_), .B(_2270_), .Q(_2038__20_) );
NO2I1X1 NO2I1X1_40 ( .gnd!(gnd!), .vdd!(vdd!), .AN(CNTR_Timer_21_), .B(_2265_), .Q(_2271_) );
NO3X1 NO3X1_10 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2263_), .B(CNTR_Timer_21_), .C(CNTR_Timer_20_), .Q(_2272_) );
ON21X1 ON21X1_293 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2271_), .B(_2272_), .C(_2195__bF_buf2), .Q(_2273_) );
NA2X1 NA2X1_621 ( .gnd!(gnd!), .vdd!(vdd!), .A(_681__21_), .B(CNTR_ld_timer_bF_buf1), .Q(_2274_) );
NA2X1 NA2X1_622 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2273_), .B(_2274_), .Q(_2038__21_) );
NO2I1X1 NO2I1X1_41 ( .gnd!(gnd!), .vdd!(vdd!), .AN(CNTR_Timer_22_), .B(_2272_), .Q(_2275_) );
NO3I1X1 NO3I1X1_2 ( .gnd!(gnd!), .vdd!(vdd!), .AN(_2055_), .B(_2263_), .C(CNTR_Timer_20_), .Q(_2276_) );
ON21X1 ON21X1_294 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2275_), .B(_2276_), .C(_2195__bF_buf2), .Q(_2277_) );
NA2X1 NA2X1_623 ( .gnd!(gnd!), .vdd!(vdd!), .A(_681__22_), .B(CNTR_ld_timer_bF_buf1), .Q(_2278_) );
NA2X1 NA2X1_624 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2277_), .B(_2278_), .Q(_2038__22_) );
INX1 INX1_168 ( .gnd!(gnd!), .vdd!(vdd!), .A(CNTR_Timer_23_), .Q(_2279_) );
AN31X1 AN31X1_70 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2266_), .B(_2055_), .C(_2267_), .D(_2279_), .Q(_2280_) );
AND4X1 AND4X1_10 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2053_), .B(_2056_), .C(_2044_), .D(_2193_), .Q(_2281_) );
ON21X1 ON21X1_295 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2280_), .B(_2281_), .C(_2195__bF_buf0), .Q(_2282_) );
NA2X1 NA2X1_625 ( .gnd!(gnd!), .vdd!(vdd!), .A(_681__23_), .B(CNTR_ld_timer_bF_buf0), .Q(_2283_) );
NA2X1 NA2X1_626 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2282_), .B(_2283_), .Q(_2038__23_) );
NO2X1 NO2X1_265 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2045_), .B(_2281_), .Q(_2284_) );
AND5X1 AND5X1_7 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2045_), .B(_2053_), .C(_2056_), .D(_2044_), .E(_2193_), .Q(_2285_) );
NO2X1 NO2X1_266 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2285_), .B(_2284_), .Q(_2286_) );
NA2X1 NA2X1_627 ( .gnd!(gnd!), .vdd!(vdd!), .A(_681__24_), .B(CNTR_ld_timer_bF_buf3), .Q(_2287_) );
ON21X1 ON21X1_296 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2286_), .B(_2192_), .C(_2287_), .Q(_2038__24_) );
INX1 INX1_169 ( .gnd!(gnd!), .vdd!(vdd!), .A(CNTR_Timer_25_), .Q(_2288_) );
NO2X1 NO2X1_267 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2288_), .B(_2285_), .Q(_2289_) );
AND2X2 AND2X2_67 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2285_), .B(_2288_), .Q(_2290_) );
ON21X1 ON21X1_297 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2290_), .B(_2289_), .C(_2195__bF_buf1), .Q(_2291_) );
NA2X1 NA2X1_628 ( .gnd!(gnd!), .vdd!(vdd!), .A(_681__25_), .B(CNTR_ld_timer_bF_buf1), .Q(_2292_) );
NA2X1 NA2X1_629 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2291_), .B(_2292_), .Q(_2038__25_) );
INX1 INX1_170 ( .gnd!(gnd!), .vdd!(vdd!), .A(CNTR_Timer_26_), .Q(_2293_) );
AN31X1 AN31X1_71 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2288_), .B(_2045_), .C(_2281_), .D(_2293_), .Q(_2294_) );
AND5X1 AND5X1_8 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2045_), .B(_2049_), .C(_2056_), .D(_2193_), .E(_2262_), .Q(_2295_) );
NO2X1 NO2X1_268 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2295_), .B(_2294_), .Q(_2296_) );
ON22X1 ON22X1_74 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2296_), .B(_2192_), .C(_2165_), .D(_2188_), .Q(_2038__26_) );
INX1 INX1_171 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2049_), .Q(_2297_) );
NA3X1 NA3X1_11 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2056_), .B(_2193_), .C(_2262_), .Q(_2298_) );
ON31X1 ON31X1_81 ( .gnd!(gnd!), .vdd!(vdd!), .A(CNTR_Timer_24_), .B(_2297_), .C(_2298_), .D(CNTR_Timer_27_), .Q(_2299_) );
NA2X1 NA2X1_630 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2295_), .B(_2046_), .Q(_2300_) );
NA2X1 NA2X1_631 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2300_), .B(_2299_), .Q(_2301_) );
NA2X1 NA2X1_632 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2301_), .B(_2195__bF_buf0), .Q(_2302_) );
NA2X1 NA2X1_633 ( .gnd!(gnd!), .vdd!(vdd!), .A(_681__27_), .B(CNTR_ld_timer_bF_buf2), .Q(_2303_) );
NA2X1 NA2X1_634 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2302_), .B(_2303_), .Q(_2038__27_) );
NO2X1 NO2X1_269 ( .gnd!(gnd!), .vdd!(vdd!), .A(CNTR_Timer_27_), .B(CNTR_Timer_28_), .Q(_2304_) );
AND3X4 AND3X4_11 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2285_), .B(_2304_), .C(_2049_), .Q(_2305_) );
INX1 INX1_172 ( .gnd!(gnd!), .vdd!(vdd!), .A(CNTR_Timer_28_), .Q(_2306_) );
AN31X1 AN31X1_72 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2046_), .B(_2049_), .C(_2285_), .D(_2306_), .Q(_2307_) );
ON21X1 ON21X1_298 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2305_), .B(_2307_), .C(_2195__bF_buf1), .Q(_2308_) );
NA2X1 NA2X1_635 ( .gnd!(gnd!), .vdd!(vdd!), .A(_681__28_), .B(CNTR_ld_timer_bF_buf1), .Q(_2309_) );
NA2X1 NA2X1_636 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2308_), .B(_2309_), .Q(_2038__28_) );
INX1 INX1_173 ( .gnd!(gnd!), .vdd!(vdd!), .A(CNTR_Timer_29_), .Q(_2310_) );
AN31X1 AN31X1_73 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2304_), .B(_2049_), .C(_2285_), .D(_2310_), .Q(_2311_) );
AND5X1 AND5X1_9 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2045_), .B(_2310_), .C(_2304_), .D(_2049_), .E(_2281_), .Q(_2312_) );
ON21X1 ON21X1_299 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2312_), .B(_2311_), .C(_2195__bF_buf1), .Q(_2313_) );
NA2X1 NA2X1_637 ( .gnd!(gnd!), .vdd!(vdd!), .A(_681__29_), .B(CNTR_ld_timer_bF_buf1), .Q(_2314_) );
NA2X1 NA2X1_638 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2313_), .B(_2314_), .Q(_2038__29_) );
INX1 INX1_174 ( .gnd!(gnd!), .vdd!(vdd!), .A(CNTR_Timer_30_), .Q(_2315_) );
AN31X1 AN31X1_74 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2310_), .B(_2304_), .C(_2295_), .D(_2315_), .Q(_2316_) );
AND5X1 AND5X1_10 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2045_), .B(_2304_), .C(_2048_), .D(_2049_), .E(_2281_), .Q(_2317_) );
ON21X1 ON21X1_300 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2316_), .B(_2317_), .C(_2195__bF_buf1), .Q(_2318_) );
NA2X1 NA2X1_639 ( .gnd!(gnd!), .vdd!(vdd!), .A(_681__30_), .B(CNTR_ld_timer_bF_buf3), .Q(_2319_) );
NA2X1 NA2X1_640 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2318_), .B(_2319_), .Q(_2038__30_) );
NA2X1 NA2X1_641 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2188_), .B(CNTR_Timer_31_), .Q(_2320_) );
ON22X1 ON22X1_75 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2317_), .B(_2320_), .C(_2185_), .D(_2188_), .Q(_2038__31_) );
INX3 INX3_8 ( .gnd!(gnd!), .vdd!(vdd!), .A(rst), .Q(_2243_) );
DFRRQX1 DFRRQX1_90 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf44), .D(_2039__0_), .Q(CNTR_gie), .RN(_2243__bF_buf7) );
DFRRQX1 DFRRQX1_91 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf7), .D(_2039__1_), .Q(CNTR_tie), .RN(_2243__bF_buf7) );
DFRRQX1 DFRRQX1_92 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf7), .D(_2039__2_), .Q(CNTR_eie), .RN(_2243__bF_buf7) );
DFRRQX1 DFRRQX1_93 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf10), .D(_2037__0_), .Q(CNTR_Cycle_0_), .RN(_2243__bF_buf7) );
DFRRQX1 DFRRQX1_94 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf17), .D(_2037__1_), .Q(CNTR_Cycle_1_), .RN(_2243__bF_buf6) );
DFRRQX1 DFRRQX1_95 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf17), .D(_2037__2_), .Q(CNTR_Cycle_2_), .RN(_2243__bF_buf6) );
DFRRQX1 DFRRQX1_96 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf6), .D(_2037__3_), .Q(CNTR_Cycle_3_), .RN(_2243__bF_buf6) );
DFRRQX1 DFRRQX1_97 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf36), .D(_2037__4_), .Q(CNTR_Cycle_4_), .RN(_2243__bF_buf4) );
DFRRQX1 DFRRQX1_98 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf36), .D(_2037__5_), .Q(CNTR_Cycle_5_), .RN(_2243__bF_buf4) );
DFRRQX1 DFRRQX1_99 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf10), .D(_2037__6_), .Q(CNTR_Cycle_6_), .RN(_2243__bF_buf7) );
DFRRQX1 DFRRQX1_100 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf36), .D(_2037__7_), .Q(CNTR_Cycle_7_), .RN(_2243__bF_buf4) );
DFRRQX1 DFRRQX1_101 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf6), .D(_2037__8_), .Q(CNTR_Cycle_8_), .RN(_2243__bF_buf6) );
DFRRQX1 DFRRQX1_102 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf6), .D(_2037__9_), .Q(CNTR_Cycle_9_), .RN(_2243__bF_buf6) );
DFRRQX1 DFRRQX1_103 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf6), .D(_2037__10_), .Q(CNTR_Cycle_10_), .RN(_2243__bF_buf6) );
DFRRQX1 DFRRQX1_104 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf47), .D(_2037__11_), .Q(CNTR_Cycle_11_), .RN(_2243__bF_buf5) );
DFRRQX1 DFRRQX1_105 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf19), .D(_2037__12_), .Q(CNTR_Cycle_12_), .RN(_2243__bF_buf5) );
DFRRQX1 DFRRQX1_106 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf19), .D(_2037__13_), .Q(CNTR_Cycle_13_), .RN(_2243__bF_buf5) );
DFRRQX1 DFRRQX1_107 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf6), .D(_2037__14_), .Q(CNTR_Cycle_14_), .RN(_2243__bF_buf1) );
DFRRQX1 DFRRQX1_108 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf19), .D(_2037__15_), .Q(CNTR_Cycle_15_), .RN(_2243__bF_buf3) );
DFRRQX1 DFRRQX1_109 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf11), .D(_2037__16_), .Q(CNTR_Cycle_16_), .RN(_2243__bF_buf1) );
DFRRQX1 DFRRQX1_110 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf47), .D(_2037__17_), .Q(CNTR_Cycle_17_), .RN(_2243__bF_buf0) );
DFRRQX1 DFRRQX1_111 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf11), .D(_2037__18_), .Q(CNTR_Cycle_18_), .RN(_2243__bF_buf1) );
DFRRQX1 DFRRQX1_112 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf47), .D(_2037__19_), .Q(CNTR_Cycle_19_), .RN(_2243__bF_buf0) );
DFRRQX1 DFRRQX1_113 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf47), .D(_2037__20_), .Q(CNTR_Cycle_20_), .RN(_2243__bF_buf0) );
DFRRQX1 DFRRQX1_114 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf47), .D(_2037__21_), .Q(CNTR_Cycle_21_), .RN(_2243__bF_buf0) );
DFRRQX1 DFRRQX1_115 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf47), .D(_2037__22_), .Q(CNTR_Cycle_22_), .RN(_2243__bF_buf0) );
DFRRQX1 DFRRQX1_116 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf11), .D(_2037__23_), .Q(CNTR_Cycle_23_), .RN(_2243__bF_buf1) );
DFRRQX1 DFRRQX1_117 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf11), .D(_2037__24_), .Q(CNTR_Cycle_24_), .RN(_2243__bF_buf1) );
DFRRQX1 DFRRQX1_118 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf6), .D(_2037__25_), .Q(CNTR_Cycle_25_), .RN(_2243__bF_buf1) );
DFRRQX1 DFRRQX1_119 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf11), .D(_2037__26_), .Q(CNTR_Cycle_26_), .RN(_2243__bF_buf1) );
DFRRQX1 DFRRQX1_120 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf17), .D(_2037__27_), .Q(CNTR_Cycle_27_), .RN(_2243__bF_buf6) );
DFRRQX1 DFRRQX1_121 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf17), .D(_2037__28_), .Q(CNTR_Cycle_28_), .RN(_2243__bF_buf1) );
DFRRQX1 DFRRQX1_122 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf6), .D(_2037__29_), .Q(CNTR_Cycle_29_), .RN(_2243__bF_buf6) );
DFRRQX1 DFRRQX1_123 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf17), .D(_2037__30_), .Q(CNTR_Cycle_30_), .RN(_2243__bF_buf6) );
DFRRQX1 DFRRQX1_124 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf19), .D(_2037__31_), .Q(CNTR_Cycle_31_), .RN(_2243__bF_buf3) );
DFRRQX1 DFRRQX1_125 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf10), .D(_2038__0_), .Q(CNTR_Timer_0_), .RN(_2243__bF_buf7) );
DFRRQX1 DFRRQX1_126 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf10), .D(_2038__1_), .Q(CNTR_Timer_1_), .RN(_2243__bF_buf7) );
DFRRQX1 DFRRQX1_127 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf10), .D(_2038__2_), .Q(CNTR_Timer_2_), .RN(_2243__bF_buf7) );
DFRRQX1 DFRRQX1_128 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf10), .D(_2038__3_), .Q(CNTR_Timer_3_), .RN(_2243__bF_buf7) );
DFRRQX1 DFRRQX1_129 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf36), .D(_2038__4_), .Q(CNTR_Timer_4_), .RN(_2243__bF_buf4) );
DFRRQX1 DFRRQX1_130 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf22), .D(_2038__5_), .Q(CNTR_Timer_5_), .RN(_2243__bF_buf4) );
DFRRQX1 DFRRQX1_131 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf22), .D(_2038__6_), .Q(CNTR_Timer_6_), .RN(_2243__bF_buf4) );
DFRRQX1 DFRRQX1_132 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf36), .D(_2038__7_), .Q(CNTR_Timer_7_), .RN(_2243__bF_buf4) );
DFRRQX1 DFRRQX1_133 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf22), .D(_2038__8_), .Q(CNTR_Timer_8_), .RN(_2243__bF_buf4) );
DFRRQX1 DFRRQX1_134 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf36), .D(_2038__9_), .Q(CNTR_Timer_9_), .RN(_2243__bF_buf3) );
DFRRQX1 DFRRQX1_135 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf36), .D(_2038__10_), .Q(CNTR_Timer_10_), .RN(_2243__bF_buf3) );
DFRRQX1 DFRRQX1_136 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf36), .D(_2038__11_), .Q(CNTR_Timer_11_), .RN(_2243__bF_buf3) );
DFRRQX1 DFRRQX1_137 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf22), .D(_2038__12_), .Q(CNTR_Timer_12_), .RN(_2243__bF_buf3) );
DFRRQX1 DFRRQX1_138 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf5), .D(_2038__13_), .Q(CNTR_Timer_13_), .RN(_2243__bF_buf2) );
DFRRQX1 DFRRQX1_139 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf22), .D(_2038__14_), .Q(CNTR_Timer_14_), .RN(_2243__bF_buf3) );
DFRRQX1 DFRRQX1_140 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf19), .D(_2038__15_), .Q(CNTR_Timer_15_), .RN(_2243__bF_buf2) );
DFRRQX1 DFRRQX1_141 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf47), .D(_2038__16_), .Q(CNTR_Timer_16_), .RN(_2243__bF_buf5) );
DFRRQX1 DFRRQX1_142 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf13), .D(_2038__17_), .Q(CNTR_Timer_17_), .RN(_2243__bF_buf0) );
DFRRQX1 DFRRQX1_143 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf13), .D(_2038__18_), .Q(CNTR_Timer_18_), .RN(_2243__bF_buf5) );
DFRRQX1 DFRRQX1_144 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf13), .D(_2038__19_), .Q(CNTR_Timer_19_), .RN(_2243__bF_buf0) );
DFRRQX1 DFRRQX1_145 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf13), .D(_2038__20_), .Q(CNTR_Timer_20_), .RN(_2243__bF_buf0) );
DFRRQX1 DFRRQX1_146 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf5), .D(_2038__21_), .Q(CNTR_Timer_21_), .RN(_2243__bF_buf2) );
DFRRQX1 DFRRQX1_147 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf5), .D(_2038__22_), .Q(CNTR_Timer_22_), .RN(_2243__bF_buf5) );
DFRRQX1 DFRRQX1_148 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf19), .D(_2038__23_), .Q(CNTR_Timer_23_), .RN(_2243__bF_buf5) );
DFRRQX1 DFRRQX1_149 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf5), .D(_2038__24_), .Q(CNTR_Timer_24_), .RN(_2243__bF_buf5) );
DFRRQX1 DFRRQX1_150 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf5), .D(_2038__25_), .Q(CNTR_Timer_25_), .RN(_2243__bF_buf2) );
DFRRQX1 DFRRQX1_151 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf19), .D(_2038__26_), .Q(CNTR_Timer_26_), .RN(_2243__bF_buf2) );
DFRRQX1 DFRRQX1_152 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf22), .D(_2038__27_), .Q(CNTR_Timer_27_), .RN(_2243__bF_buf2) );
DFRRQX1 DFRRQX1_153 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf5), .D(_2038__28_), .Q(CNTR_Timer_28_), .RN(_2243__bF_buf2) );
DFRRQX1 DFRRQX1_154 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf5), .D(_2038__29_), .Q(CNTR_Timer_29_), .RN(_2243__bF_buf2) );
DFRRQX1 DFRRQX1_155 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf47), .D(_2038__30_), .Q(CNTR_Timer_30_), .RN(_2243__bF_buf5) );
DFRRQX1 DFRRQX1_156 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf22), .D(_2038__31_), .Q(CNTR_Timer_31_), .RN(_2243__bF_buf3) );
NO2X1 NO2X1_270 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_IDEC0_IR_2_), .B(_686__0_), .Q(_2330_) );
NO2X1 NO2X1_271 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_IDEC0_IR_7_), .B(CTRL_IDEC0_IR_3_), .Q(_2331_) );
NO2X1 NO2X1_272 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_IDEC0_IR_8_), .B(CTRL_IDEC0_IR_11_), .Q(_2332_) );
NO2X1 NO2X1_273 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_IDEC0_IR_9_), .B(CTRL_IDEC0_IR_10_), .Q(_2333_) );
AND4X1 AND4X1_11 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2330_), .B(_2331_), .C(_2332_), .D(_2333_), .Q(_2334_) );
NO2X1 NO2X1_274 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_IDEC0_IR_13_), .B(CTRL_IDEC0_IR_12_), .Q(_2335_) );
NA3I1X1 NA3I1X1_101 ( .gnd!(gnd!), .vdd!(vdd!), .AN(CTRL_IDEC0_IR_14_), .B(CTRL_IDEC0_IR_0_), .C(_2335_), .Q(_2336_) );
AND4X1 AND4X1_12 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_IDEC0_IR_4_), .B(CTRL_IDEC0_IR_1_), .C(CTRL_IDEC0_IR_6_), .D(CTRL_IDEC0_IR_5_), .Q(_2337_) );
NA3I1X1 NA3I1X1_102 ( .gnd!(gnd!), .vdd!(vdd!), .AN(_2336_), .B(_2337_), .C(_2334_), .Q(_2338_) );
NO2X1 NO2X1_275 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_IDEC0_IR_25_), .B(_687__4_), .Q(_2339_) );
NO2X1 NO2X1_276 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_IDEC0_IR_27_), .B(CTRL_IDEC0_IR_26_), .Q(_2340_) );
NO2X1 NO2X1_277 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_IDEC0_IR_28_), .B(CTRL_IDEC0_IR_31_), .Q(_2341_) );
NO2X1 NO2X1_278 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_IDEC0_IR_29_), .B(CTRL_IDEC0_IR_30_), .Q(_2342_) );
AND4X1 AND4X1_13 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2339_), .B(_2340_), .C(_2341_), .D(_2342_), .Q(_2343_) );
NO2X1 NO2X1_279 ( .gnd!(gnd!), .vdd!(vdd!), .A(_686__1_), .B(_686__4_), .Q(_2344_) );
NO2X1 NO2X1_280 ( .gnd!(gnd!), .vdd!(vdd!), .A(_686__2_), .B(_686__3_), .Q(_2345_) );
AND2X2 AND2X2_68 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2344_), .B(_2345_), .Q(_2346_) );
NO2X1 NO2X1_281 ( .gnd!(gnd!), .vdd!(vdd!), .A(_687__3_), .B(_687__2_), .Q(_2347_) );
NA3I1X1 NA3I1X1_103 ( .gnd!(gnd!), .vdd!(vdd!), .AN(_687__0_), .B(_687__1_), .C(_2347_), .Q(_2348_) );
NA3I1X1 NA3I1X1_104 ( .gnd!(gnd!), .vdd!(vdd!), .AN(_2348_), .B(_2346_), .C(_2343_), .Q(_2349_) );
NO2X2 NO2X2_3 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2338_), .B(_2349_), .Q(CTRL_cu_pc_s4) );
NO2X1 NO2X1_282 ( .gnd!(gnd!), .vdd!(vdd!), .A(_687__0_), .B(_687__1_), .Q(_2350_) );
AND4X1 AND4X1_14 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2344_), .B(_2345_), .C(_2347_), .D(_2350_), .Q(_2351_) );
NA2X1 NA2X1_642 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2343_), .B(_2351_), .Q(_2352_) );
NO2X1 NO2X1_283 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2352_), .B(_2338_), .Q(CTRL_cu_int_ecall) );
NA2X1 NA2X1_643 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2344_), .B(_2345_), .Q(_2353_) );
NA3I1X1 NA3I1X1_105 ( .gnd!(gnd!), .vdd!(vdd!), .AN(_687__1_), .B(_687__0_), .C(_2347_), .Q(_2354_) );
NO2X1 NO2X1_284 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2353_), .B(_2354_), .Q(_2355_) );
NA2X1 NA2X1_644 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2355_), .B(_2343_), .Q(_2356_) );
NO2X1 NO2X1_285 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2356_), .B(_2338_), .Q(CTRL_cu_int_ebreak) );
INX2 INX2_11 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_cyc_bF_buf7_bF_buf2), .Q(_2329_) );
ON31X1 ON31X1_82 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_IDEC1_cu_alu_i_inst), .B(CTRL_IDEC1_cu_alu_r_inst), .C(CTRL_IDEC1_cu_br_inst), .D(_2329__bF_buf3), .Q(_2357_) );
MU2X1 MU2X1_205 ( .gnd!(gnd!), .vdd!(vdd!), .IN0(ALU_cf), .IN1(CTRL_BR_cf), .Q(_2321_), .S(_2357_) );
MU2X1 MU2X1_206 ( .gnd!(gnd!), .vdd!(vdd!), .IN0(ALU_sf), .IN1(CTRL_BR_sf), .Q(_2325_), .S(_2357_) );
MU2X1 MU2X1_207 ( .gnd!(gnd!), .vdd!(vdd!), .IN0(ALU_zf), .IN1(CTRL_BR_zf), .Q(_2328_), .S(_2357_) );
MU2X1 MU2X1_208 ( .gnd!(gnd!), .vdd!(vdd!), .IN0(ALU_vf), .IN1(CTRL_BR_vf), .Q(_2327_), .S(_2357_) );
MU2X1 MU2X1_209 ( .gnd!(gnd!), .vdd!(vdd!), .IN0(CTRL_IDEC2_IR_2_), .IN1(ALU_opcode_0_), .Q(_2323__2_), .S(CTRL_cyc_bF_buf6_bF_buf3) );
MU2X1 MU2X1_210 ( .gnd!(gnd!), .vdd!(vdd!), .IN0(CTRL_IDEC2_IR_3_), .IN1(ALU_opcode_1_), .Q(_2323__3_), .S(CTRL_cyc_bF_buf5_bF_buf1) );
MU2X1 MU2X1_211 ( .gnd!(gnd!), .vdd!(vdd!), .IN0(CTRL_IDEC2_IR_4_), .IN1(ALU_opcode_2_), .Q(_2323__4_), .S(CTRL_cyc_bF_buf4_bF_buf2) );
MU2X1 MU2X1_212 ( .gnd!(gnd!), .vdd!(vdd!), .IN0(CTRL_IDEC2_IR_5_), .IN1(ALU_opcode_3_), .Q(_2323__5_), .S(CTRL_cyc_bF_buf3_bF_buf0) );
MU2X1 MU2X1_213 ( .gnd!(gnd!), .vdd!(vdd!), .IN0(CTRL_IDEC2_IR_6_), .IN1(ALU_opcode_4_), .Q(_2323__6_), .S(CTRL_cyc_bF_buf2_bF_buf3) );
MU2X1 MU2X1_214 ( .gnd!(gnd!), .vdd!(vdd!), .IN0(_685__0_), .IN1(CTRL_IDEC1_IR_7_), .Q(_2323__7_), .S(CTRL_cyc_bF_buf1_bF_buf3) );
MU2X1 MU2X1_215 ( .gnd!(gnd!), .vdd!(vdd!), .IN0(_685__1_), .IN1(CTRL_IDEC1_IR_8_), .Q(_2323__8_), .S(CTRL_cyc_bF_buf0_bF_buf0) );
INX1 INX1_175 ( .gnd!(gnd!), .vdd!(vdd!), .A(_685__2_), .Q(_2358_) );
INX1 INX1_176 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_IDEC1_IR_9_), .Q(_2359_) );
MU2IX1 MU2IX1_108 ( .gnd!(gnd!), .vdd!(vdd!), .IN0(_2358_), .IN1(_2359_), .Q(_2323__9_), .S(CTRL_cyc_bF_buf14_bF_buf2) );
MU2X1 MU2X1_216 ( .gnd!(gnd!), .vdd!(vdd!), .IN0(_685__3_), .IN1(CTRL_IDEC1_IR_10_), .Q(_2323__10_), .S(CTRL_cyc_bF_buf13_bF_buf3) );
INX1 INX1_177 ( .gnd!(gnd!), .vdd!(vdd!), .A(_685__4_), .Q(_2360_) );
INX1 INX1_178 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_IDEC1_IR_11_), .Q(_2361_) );
MU2IX1 MU2IX1_109 ( .gnd!(gnd!), .vdd!(vdd!), .IN0(_2360_), .IN1(_2361_), .Q(_2323__11_), .S(CTRL_cyc_bF_buf12_bF_buf3) );
INX1 INX1_179 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_IDEC1_cu_custom_inst_bF_buf3), .Q(_2362_) );
NO2X3 NO2X3_1 ( .gnd!(gnd!), .vdd!(vdd!), .A(extDone), .B(_2362_), .Q(CTRL_cu_ext_hold) );
AN22X1 AN22X1_69 ( .gnd!(gnd!), .vdd!(vdd!), .A(CNTR_tie), .B(CTRL_TMRIF), .C(CNTR_eie), .D(IRQ), .Q(_2363_) );
ON21X1 ON21X1_301 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2355_), .B(_2351_), .C(_2343_), .Q(_2364_) );
ON21X1 ON21X1_302 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2364_), .B(_2338_), .C(_2363_), .Q(_2365_) );
NO2I1X1 NO2I1X1_42 ( .gnd!(gnd!), .vdd!(vdd!), .AN(CNTR_gie), .B(CTRL_ISRMode), .Q(_2366_) );
NA2X2 NA2X2_3 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2365_), .B(_2366_), .Q(_2367_) );
INX1 INX1_180 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2367__bF_buf2), .Q(CTRL_cu_pc_s0) );
INX1 INX1_181 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_IDEC1_cu_jal_inst), .Q(_2368_) );
NA2I1X1 NA2I1X1_80 ( .gnd!(gnd!), .vdd!(vdd!), .AN(CTRL_IDEC1_cu_jalr_inst_bF_buf4), .B(_2368_), .Q(CTRL_cu_j_inst_1) );
NO2X1 NO2X1_286 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_IDEC1_cu_br_inst), .B(CTRL_cu_j_inst_1), .Q(_2369_) );
NA2X1 NA2X1_645 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2329__bF_buf2), .B(ALU_opcode_0_), .Q(_2370_) );
INX1 INX1_182 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2369_), .Q(_2371_) );
NA2I1X1 NA2I1X1_81 ( .gnd!(gnd!), .vdd!(vdd!), .AN(ALU_opcode_0_), .B(CTRL_cu_ext_hold_bF_buf6), .Q(_2372_) );
ON211X1 ON211X1_84 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_IDEC0_IR_2_), .B(CTRL_cu_ext_hold_bF_buf6), .C(_2372_), .D(CTRL_cyc_bF_buf11_bF_buf1), .Q(_2373_) );
NA3I2X1 NA3I2X1_2 ( .gnd!(gnd!), .vdd!(vdd!), .AN(_2371__bF_buf1), .BN(_2373_), .C(_2367__bF_buf3), .Q(_2374_) );
NA2X1 NA2X1_646 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2374_), .B(_2370_), .Q(_2322__2_) );
NA2X1 NA2X1_647 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2329__bF_buf3), .B(ALU_opcode_1_), .Q(_2375_) );
NA2I1X1 NA2I1X1_82 ( .gnd!(gnd!), .vdd!(vdd!), .AN(ALU_opcode_1_), .B(CTRL_cu_ext_hold_bF_buf2), .Q(_2376_) );
ON211X1 ON211X1_85 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_IDEC0_IR_3_), .B(CTRL_cu_ext_hold_bF_buf2), .C(_2376_), .D(CTRL_cyc_bF_buf10_bF_buf0), .Q(_2377_) );
NA3I2X1 NA3I2X1_3 ( .gnd!(gnd!), .vdd!(vdd!), .AN(_2371__bF_buf3), .BN(_2377_), .C(_2367__bF_buf2), .Q(_2378_) );
NA2X1 NA2X1_648 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2378_), .B(_2375_), .Q(_2322__3_) );
MU2X1 MU2X1_217 ( .gnd!(gnd!), .vdd!(vdd!), .IN0(CTRL_IDEC0_IR_4_), .IN1(ALU_opcode_2_), .Q(_2379_), .S(CTRL_cu_ext_hold_bF_buf5) );
NO2X1 NO2X1_287 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2329__bF_buf3), .B(_2379_), .Q(_2380_) );
NO2X1 NO2X1_288 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_cyc_bF_buf9_bF_buf3), .B(ALU_opcode_2_), .Q(_2381_) );
AN31X1 AN31X1_75 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2369_), .B(_2380_), .C(_2367__bF_buf0), .D(_2381_), .Q(_2322__4_) );
NA2X1 NA2X1_649 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2329__bF_buf2), .B(ALU_opcode_3_), .Q(_2382_) );
NA2I1X1 NA2I1X1_83 ( .gnd!(gnd!), .vdd!(vdd!), .AN(ALU_opcode_3_), .B(CTRL_cu_ext_hold_bF_buf1), .Q(_2383_) );
ON211X1 ON211X1_86 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_IDEC0_IR_5_), .B(CTRL_cu_ext_hold_bF_buf5), .C(_2383_), .D(CTRL_cyc_bF_buf8_bF_buf3), .Q(_2384_) );
NA3I2X1 NA3I2X1_4 ( .gnd!(gnd!), .vdd!(vdd!), .AN(_2371__bF_buf1), .BN(_2384_), .C(_2367__bF_buf3), .Q(_2385_) );
NA2X1 NA2X1_650 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2385_), .B(_2382_), .Q(_2322__5_) );
NA2X1 NA2X1_651 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2329__bF_buf2), .B(ALU_opcode_4_), .Q(_2386_) );
NA2I1X1 NA2I1X1_84 ( .gnd!(gnd!), .vdd!(vdd!), .AN(ALU_opcode_4_), .B(CTRL_cu_ext_hold_bF_buf6), .Q(_2387_) );
ON211X1 ON211X1_87 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_IDEC0_IR_6_), .B(CTRL_cu_ext_hold_bF_buf6), .C(_2387_), .D(CTRL_cyc_bF_buf7_bF_buf2), .Q(_2388_) );
NA3I2X1 NA3I2X1_5 ( .gnd!(gnd!), .vdd!(vdd!), .AN(_2371__bF_buf1), .BN(_2388_), .C(_2367__bF_buf3), .Q(_2389_) );
NA2X1 NA2X1_652 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2389_), .B(_2386_), .Q(_2322__6_) );
NA2X1 NA2X1_653 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2329__bF_buf4), .B(CTRL_IDEC1_IR_7_), .Q(_2390_) );
INX1 INX1_183 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_IDEC1_IR_7_), .Q(_2391_) );
NA2X1 NA2X1_654 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_cu_ext_hold_bF_buf0), .B(_2391_), .Q(_2392_) );
ON211X1 ON211X1_88 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_IDEC0_IR_7_), .B(CTRL_cu_ext_hold_bF_buf3), .C(_2392_), .D(CTRL_cyc_bF_buf6_bF_buf3), .Q(_2393_) );
NA3I2X1 NA3I2X1_6 ( .gnd!(gnd!), .vdd!(vdd!), .AN(_2371__bF_buf2), .BN(_2393_), .C(_2367__bF_buf1), .Q(_2394_) );
NA2X1 NA2X1_655 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2394_), .B(_2390_), .Q(_2322__7_) );
NA2X1 NA2X1_656 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2329__bF_buf4), .B(CTRL_IDEC1_IR_8_), .Q(_2395_) );
NA2I1X1 NA2I1X1_85 ( .gnd!(gnd!), .vdd!(vdd!), .AN(CTRL_IDEC1_IR_8_), .B(CTRL_cu_ext_hold_bF_buf3), .Q(_2396_) );
ON211X1 ON211X1_89 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_IDEC0_IR_8_), .B(CTRL_cu_ext_hold_bF_buf1), .C(_2396_), .D(CTRL_cyc_bF_buf5_bF_buf3), .Q(_2397_) );
NA3I2X1 NA3I2X1_7 ( .gnd!(gnd!), .vdd!(vdd!), .AN(_2371__bF_buf2), .BN(_2397_), .C(_2367__bF_buf1), .Q(_2398_) );
NA2X1 NA2X1_657 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2398_), .B(_2395_), .Q(_2322__8_) );
NA2X1 NA2X1_658 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2329__bF_buf4), .B(CTRL_IDEC1_IR_9_), .Q(_2399_) );
NA2X1 NA2X1_659 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_cu_ext_hold_bF_buf0), .B(_2359_), .Q(_2400_) );
ON211X1 ON211X1_90 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_IDEC0_IR_9_), .B(CTRL_cu_ext_hold_bF_buf0), .C(_2400_), .D(CTRL_cyc_bF_buf4_bF_buf2), .Q(_2401_) );
NA3I2X1 NA3I2X1_8 ( .gnd!(gnd!), .vdd!(vdd!), .AN(_2371__bF_buf0), .BN(_2401_), .C(_2367__bF_buf4), .Q(_2402_) );
NA2X1 NA2X1_660 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2402_), .B(_2399_), .Q(_2322__9_) );
NA2X1 NA2X1_661 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2329__bF_buf2), .B(CTRL_IDEC1_IR_10_), .Q(_2403_) );
NA2I1X1 NA2I1X1_86 ( .gnd!(gnd!), .vdd!(vdd!), .AN(CTRL_IDEC1_IR_10_), .B(CTRL_cu_ext_hold_bF_buf4), .Q(_2404_) );
ON211X1 ON211X1_91 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_IDEC0_IR_10_), .B(CTRL_cu_ext_hold_bF_buf4), .C(_2404_), .D(CTRL_cyc_bF_buf3_bF_buf0), .Q(_2405_) );
NA3I2X1 NA3I2X1_9 ( .gnd!(gnd!), .vdd!(vdd!), .AN(_2371__bF_buf2), .BN(_2405_), .C(_2367__bF_buf1), .Q(_2406_) );
NA2X1 NA2X1_662 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2406_), .B(_2403_), .Q(_2322__10_) );
NA2X1 NA2X1_663 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2329__bF_buf1), .B(CTRL_IDEC1_IR_11_), .Q(_2407_) );
NA2X1 NA2X1_664 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_cu_ext_hold_bF_buf4), .B(_2361_), .Q(_2408_) );
ON211X1 ON211X1_92 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_IDEC0_IR_11_), .B(CTRL_cu_ext_hold_bF_buf4), .C(_2408_), .D(CTRL_cyc_bF_buf2_bF_buf3), .Q(_2409_) );
NA3I2X1 NA3I2X1_10 ( .gnd!(gnd!), .vdd!(vdd!), .AN(_2371__bF_buf1), .BN(_2409_), .C(_2367__bF_buf3), .Q(_2410_) );
NA2X1 NA2X1_665 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2410_), .B(_2407_), .Q(_2322__11_) );
NA2X1 NA2X1_666 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2329__bF_buf0), .B(_682__0_bF_buf3), .Q(_2411_) );
NA2I1X1 NA2I1X1_87 ( .gnd!(gnd!), .vdd!(vdd!), .AN(_682__0_bF_buf3), .B(CTRL_cu_ext_hold_bF_buf5), .Q(_2412_) );
ON211X1 ON211X1_93 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_IDEC0_IR_12_), .B(CTRL_cu_ext_hold_bF_buf1), .C(_2412_), .D(CTRL_cyc_bF_buf1_bF_buf3), .Q(_2413_) );
NA3I2X1 NA3I2X1_11 ( .gnd!(gnd!), .vdd!(vdd!), .AN(_2371__bF_buf0), .BN(_2413_), .C(_2367__bF_buf0), .Q(_2414_) );
NA2X1 NA2X1_667 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2414_), .B(_2411_), .Q(_2322__12_) );
NA2X1 NA2X1_668 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2329__bF_buf0), .B(_682__1_bF_buf2), .Q(_2415_) );
INX1 INX1_184 ( .gnd!(gnd!), .vdd!(vdd!), .A(_682__1_bF_buf2), .Q(_2416_) );
NA2X1 NA2X1_669 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_cu_ext_hold_bF_buf6), .B(_2416_), .Q(_2417_) );
ON211X1 ON211X1_94 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_IDEC0_IR_13_), .B(CTRL_cu_ext_hold_bF_buf2), .C(_2417_), .D(CTRL_cyc_bF_buf0_bF_buf0), .Q(_2418_) );
NA3I2X1 NA3I2X1_12 ( .gnd!(gnd!), .vdd!(vdd!), .AN(_2371__bF_buf3), .BN(_2418_), .C(_2367__bF_buf0), .Q(_2419_) );
NA2X1 NA2X1_670 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2419_), .B(_2415_), .Q(_2322__13_) );
NA2X1 NA2X1_671 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2329__bF_buf0), .B(EXT_type_bF_buf0), .Q(_2420_) );
INX1 INX1_185 ( .gnd!(gnd!), .vdd!(vdd!), .A(EXT_type_bF_buf0), .Q(_2421_) );
NA2X1 NA2X1_672 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_cu_ext_hold_bF_buf5), .B(_2421_), .Q(_2422_) );
ON211X1 ON211X1_95 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_IDEC0_IR_14_), .B(CTRL_cu_ext_hold_bF_buf5), .C(_2422_), .D(CTRL_cyc_bF_buf14_bF_buf1), .Q(_2423_) );
NA3I2X1 NA3I2X1_13 ( .gnd!(gnd!), .vdd!(vdd!), .AN(_2371__bF_buf3), .BN(_2423_), .C(_2367__bF_buf0), .Q(_2424_) );
NA2X1 NA2X1_673 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2424_), .B(_2420_), .Q(_2322__14_) );
NA2X1 NA2X1_674 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2329__bF_buf3), .B(CTRL_cu_csr_rd_s1_bF_buf2), .Q(_2425_) );
NA2I1X1 NA2I1X1_88 ( .gnd!(gnd!), .vdd!(vdd!), .AN(CTRL_cu_csr_rd_s1_bF_buf2), .B(CTRL_cu_ext_hold_bF_buf1), .Q(_2426_) );
ON211X1 ON211X1_96 ( .gnd!(gnd!), .vdd!(vdd!), .A(_687__0_), .B(CTRL_cu_ext_hold_bF_buf1), .C(_2426_), .D(CTRL_cyc_bF_buf13_bF_buf3), .Q(_2427_) );
NA3I2X1 NA3I2X1_14 ( .gnd!(gnd!), .vdd!(vdd!), .AN(_2371__bF_buf0), .BN(_2427_), .C(_2367__bF_buf4), .Q(_2428_) );
NA2X1 NA2X1_675 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2428_), .B(_2425_), .Q(_2322__20_) );
NA2X1 NA2X1_676 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2329__bF_buf1), .B(ALU_shamt_1_), .Q(_2429_) );
INX1 INX1_186 ( .gnd!(gnd!), .vdd!(vdd!), .A(ALU_shamt_1_), .Q(_2430_) );
NA2X1 NA2X1_677 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_cu_ext_hold_bF_buf3), .B(_2430_), .Q(_2431_) );
ON211X1 ON211X1_97 ( .gnd!(gnd!), .vdd!(vdd!), .A(_687__1_), .B(CTRL_cu_ext_hold_bF_buf3), .C(_2431_), .D(CTRL_cyc_bF_buf12_bF_buf3), .Q(_2432_) );
NA3I2X1 NA3I2X1_15 ( .gnd!(gnd!), .vdd!(vdd!), .AN(_2371__bF_buf2), .BN(_2432_), .C(_2367__bF_buf1), .Q(_2433_) );
NA2X1 NA2X1_678 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2433_), .B(_2429_), .Q(_2322__21_) );
NA2X1 NA2X1_679 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2329__bF_buf4), .B(ALU_shamt_2_), .Q(_2434_) );
NA2I1X1 NA2I1X1_89 ( .gnd!(gnd!), .vdd!(vdd!), .AN(ALU_shamt_2_), .B(CTRL_cu_ext_hold_bF_buf3), .Q(_2435_) );
ON211X1 ON211X1_98 ( .gnd!(gnd!), .vdd!(vdd!), .A(_687__2_), .B(CTRL_cu_ext_hold_bF_buf0), .C(_2435_), .D(CTRL_cyc_bF_buf11_bF_buf1), .Q(_2436_) );
NA3I2X1 NA3I2X1_16 ( .gnd!(gnd!), .vdd!(vdd!), .AN(_2371__bF_buf2), .BN(_2436_), .C(_2367__bF_buf4), .Q(_2437_) );
NA2X1 NA2X1_680 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2437_), .B(_2434_), .Q(_2322__22_) );
NA2X1 NA2X1_681 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2329__bF_buf0), .B(ALU_shamt_3_), .Q(_2438_) );
NA2I1X1 NA2I1X1_90 ( .gnd!(gnd!), .vdd!(vdd!), .AN(ALU_shamt_3_), .B(CTRL_cu_ext_hold_bF_buf2), .Q(_2439_) );
ON211X1 ON211X1_99 ( .gnd!(gnd!), .vdd!(vdd!), .A(_687__3_), .B(CTRL_cu_ext_hold_bF_buf2), .C(_2439_), .D(CTRL_cyc_bF_buf10_bF_buf0), .Q(_2440_) );
NA3I2X1 NA3I2X1_17 ( .gnd!(gnd!), .vdd!(vdd!), .AN(_2371__bF_buf3), .BN(_2440_), .C(_2367__bF_buf2), .Q(_2441_) );
NA2X1 NA2X1_682 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2441_), .B(_2438_), .Q(_2322__23_) );
NA2X1 NA2X1_683 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2329__bF_buf0), .B(ALU_shamt_4_), .Q(_2442_) );
NA2I1X1 NA2I1X1_91 ( .gnd!(gnd!), .vdd!(vdd!), .AN(ALU_shamt_4_), .B(CTRL_cu_ext_hold_bF_buf2), .Q(_2443_) );
ON211X1 ON211X1_100 ( .gnd!(gnd!), .vdd!(vdd!), .A(_687__4_), .B(CTRL_cu_ext_hold_bF_buf5), .C(_2443_), .D(CTRL_cyc_bF_buf9_bF_buf3), .Q(_2444_) );
NA3I2X1 NA3I2X1_18 ( .gnd!(gnd!), .vdd!(vdd!), .AN(_2371__bF_buf3), .BN(_2444_), .C(_2367__bF_buf0), .Q(_2445_) );
NA2X1 NA2X1_684 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2445_), .B(_2442_), .Q(_2322__24_) );
NA2X1 NA2X1_685 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2329__bF_buf1), .B(ALU_func7_0_), .Q(_2446_) );
NA2I1X1 NA2I1X1_92 ( .gnd!(gnd!), .vdd!(vdd!), .AN(ALU_func7_0_), .B(CTRL_cu_ext_hold_bF_buf5), .Q(_2447_) );
ON211X1 ON211X1_101 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_IDEC0_IR_25_), .B(CTRL_cu_ext_hold_bF_buf5), .C(_2447_), .D(CTRL_cyc_bF_buf8_bF_buf3), .Q(_2448_) );
NA3I2X1 NA3I2X1_19 ( .gnd!(gnd!), .vdd!(vdd!), .AN(_2371__bF_buf1), .BN(_2448_), .C(_2367__bF_buf2), .Q(_2449_) );
NA2X1 NA2X1_686 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2449_), .B(_2446_), .Q(_2322__25_) );
NA2X1 NA2X1_687 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2329__bF_buf1), .B(ALU_func7_1_), .Q(_2450_) );
NA2I1X1 NA2I1X1_93 ( .gnd!(gnd!), .vdd!(vdd!), .AN(ALU_func7_1_), .B(CTRL_cu_ext_hold_bF_buf4), .Q(_2451_) );
ON211X1 ON211X1_102 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_IDEC0_IR_26_), .B(CTRL_cu_ext_hold_bF_buf4), .C(_2451_), .D(CTRL_cyc_bF_buf7_bF_buf2), .Q(_2452_) );
NA3I2X1 NA3I2X1_20 ( .gnd!(gnd!), .vdd!(vdd!), .AN(_2371__bF_buf1), .BN(_2452_), .C(_2367__bF_buf3), .Q(_2453_) );
NA2X1 NA2X1_688 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2453_), .B(_2450_), .Q(_2322__26_) );
NA2X1 NA2X1_689 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2329__bF_buf1), .B(CTRL_cu_csr_rd_s2), .Q(_2454_) );
NA2I1X1 NA2I1X1_94 ( .gnd!(gnd!), .vdd!(vdd!), .AN(CTRL_cu_csr_rd_s2), .B(CTRL_cu_ext_hold_bF_buf6), .Q(_2455_) );
ON211X1 ON211X1_103 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_IDEC0_IR_27_), .B(CTRL_cu_ext_hold_bF_buf3), .C(_2455_), .D(CTRL_cyc_bF_buf6_bF_buf3), .Q(_2456_) );
NA3I2X1 NA3I2X1_21 ( .gnd!(gnd!), .vdd!(vdd!), .AN(_2371__bF_buf2), .BN(_2456_), .C(_2367__bF_buf1), .Q(_2457_) );
NA2X1 NA2X1_690 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2457_), .B(_2454_), .Q(_2322__27_) );
NA2X1 NA2X1_691 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2329__bF_buf4), .B(ALU_func7_3_), .Q(_2459_) );
NA2I1X1 NA2I1X1_95 ( .gnd!(gnd!), .vdd!(vdd!), .AN(ALU_func7_3_), .B(CTRL_cu_ext_hold_bF_buf3), .Q(_2460_) );
ON211X1 ON211X1_104 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_IDEC0_IR_28_), .B(CTRL_cu_ext_hold_bF_buf1), .C(_2460_), .D(CTRL_cyc_bF_buf5_bF_buf3), .Q(_2461_) );
NA3I2X1 NA3I2X1_22 ( .gnd!(gnd!), .vdd!(vdd!), .AN(_2371__bF_buf0), .BN(_2461_), .C(_2367__bF_buf4), .Q(_2462_) );
NA2X1 NA2X1_692 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2462_), .B(_2459_), .Q(_2322__28_) );
NA2X1 NA2X1_693 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2329__bF_buf4), .B(ALU_func7_4_), .Q(_2463_) );
NA2I1X1 NA2I1X1_96 ( .gnd!(gnd!), .vdd!(vdd!), .AN(ALU_func7_4_), .B(CTRL_cu_ext_hold_bF_buf0), .Q(_2464_) );
ON211X1 ON211X1_105 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_IDEC0_IR_29_), .B(CTRL_cu_ext_hold_bF_buf1), .C(_2464_), .D(CTRL_cyc_bF_buf4_bF_buf2), .Q(_2465_) );
NA3I2X1 NA3I2X1_23 ( .gnd!(gnd!), .vdd!(vdd!), .AN(_2371__bF_buf0), .BN(_2465_), .C(_2367__bF_buf4), .Q(_2466_) );
NA2X1 NA2X1_694 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2466_), .B(_2463_), .Q(_2322__29_) );
NA2X1 NA2X1_695 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2329__bF_buf1), .B(ALU_func7_5_bF_buf3), .Q(_2467_) );
NA2I1X1 NA2I1X1_97 ( .gnd!(gnd!), .vdd!(vdd!), .AN(ALU_func7_5_bF_buf3), .B(CTRL_cu_ext_hold_bF_buf6), .Q(_2468_) );
ON211X1 ON211X1_106 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_IDEC0_IR_30_), .B(CTRL_cu_ext_hold_bF_buf2), .C(_2468_), .D(CTRL_cyc_bF_buf3_bF_buf0), .Q(_2469_) );
NA3I2X1 NA3I2X1_24 ( .gnd!(gnd!), .vdd!(vdd!), .AN(_2371__bF_buf3), .BN(_2469_), .C(_2367__bF_buf2), .Q(_2470_) );
NA2X1 NA2X1_696 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2470_), .B(_2467_), .Q(_2322__30_) );
NA2X1 NA2X1_697 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2329__bF_buf4), .B(ALU_func7_6_), .Q(_2471_) );
NA2I1X1 NA2I1X1_98 ( .gnd!(gnd!), .vdd!(vdd!), .AN(ALU_func7_6_), .B(CTRL_cu_ext_hold_bF_buf0), .Q(_2472_) );
ON211X1 ON211X1_107 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_IDEC0_IR_31_), .B(CTRL_cu_ext_hold_bF_buf0), .C(_2472_), .D(CTRL_cyc_bF_buf2_bF_buf3), .Q(_2473_) );
NA3I2X1 NA3I2X1_25 ( .gnd!(gnd!), .vdd!(vdd!), .AN(_2371__bF_buf0), .BN(_2473_), .C(_2367__bF_buf4), .Q(_2474_) );
NA2X1 NA2X1_698 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2474_), .B(_2471_), .Q(_2322__31_) );
NA3I1X1 NA3I1X1_106 ( .gnd!(gnd!), .vdd!(vdd!), .AN(_2329__bF_buf0), .B(_2366_), .C(_2365_), .Q(_2475_) );
NA2I1X1 NA2I1X1_99 ( .gnd!(gnd!), .vdd!(vdd!), .AN(CTRL_cu_pc_s4_bF_buf2), .B(CTRL_ISRMode), .Q(_2476_) );
AN21X1 AN21X1_150 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2476_), .B(_2475_), .C(rst), .Q(_2324_) );
INX1 INX1_187 ( .gnd!(gnd!), .vdd!(vdd!), .A(CNTR_tif), .Q(_2477_) );
NO2X1 NO2X1_289 ( .gnd!(gnd!), .vdd!(vdd!), .A(ALU_func7_1_), .B(CTRL_cu_csr_rd_s2), .Q(_2478_) );
NO2X1 NO2X1_290 ( .gnd!(gnd!), .vdd!(vdd!), .A(ALU_shamt_4_), .B(ALU_func7_0_), .Q(_2479_) );
AND4X1 AND4X1_15 ( .gnd!(gnd!), .vdd!(vdd!), .A(_682__0_bF_buf3), .B(CTRL_IDEC1_cu_system_inst_bF_buf3), .C(_2416_), .D(_2421_), .Q(_2480_) );
NA3X1 NA3X1_12 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2478_), .B(_2479_), .C(_2480_), .Q(_2481_) );
NO2X1 NO2X1_291 ( .gnd!(gnd!), .vdd!(vdd!), .A(ALU_func7_3_), .B(ALU_func7_4_), .Q(_2482_) );
AND3X4 AND3X4_12 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2482_), .B(ALU_func7_5_bF_buf3), .C(ALU_func7_6_), .Q(_2483_) );
NO2X1 NO2X1_292 ( .gnd!(gnd!), .vdd!(vdd!), .A(ALU_shamt_2_), .B(ALU_shamt_3_), .Q(_2484_) );
AND3X4 AND3X4_13 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2430_), .B(CTRL_cu_csr_rd_s1_bF_buf2), .C(_2484_), .Q(_2485_) );
NA2X1 NA2X1_699 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2485_), .B(_2483_), .Q(_2486_) );
ON31X1 ON31X1_83 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2329__bF_buf3), .B(_2486_), .C(_2481_), .D(CTRL_TMRIF), .Q(_2487_) );
AN21X1 AN21X1_151 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2487_), .B(_2477_), .C(rst), .Q(_2326_) );
AND2X2 AND2X2_69 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_cyc_bF_buf1_bF_buf2), .B(CTRL_IDEC1_cu_store_inst), .Q(_680_) );
OR2X2 OR2X2_16 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_cu_int_ecall), .B(CTRL_cu_int_ebreak), .Q(CTRL_cu_sel_epc) );
NO2X1 NO2X1_293 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2486_), .B(_2481_), .Q(CNTR_ld_timer) );
NA2X1 NA2X1_700 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_IDEC1_cu_br_inst), .B(CTRL_BR_taken), .Q(_2488_) );
NA2X3 NA2X3_4 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2368_), .B(_2488_), .Q(CTRL_cu_pc_s2) );
NO2I1X2 NO2I1X2_1 ( .gnd!(gnd!), .vdd!(vdd!), .AN(CTRL_IDEC1_cu_br_inst), .B(CTRL_BR_taken), .Q(CTRL_cu_pc_s3) );
OR2X2 OR2X2_17 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_IDEC2_cu_alu_i_inst), .B(CTRL_IDEC2_cu_alu_r_inst), .Q(_2489_) );
NO3X1 NO3X1_11 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2489_), .B(CTRL_IDEC2_cu_jalr_inst), .C(CTRL_IDEC2_cu_jal_inst), .Q(_2490_) );
NO2X1 NO2X1_294 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_IDEC2_cu_load_inst), .B(CTRL_IDEC2_cu_auipc_inst), .Q(_2491_) );
AN211X1 AN211X1_13 ( .gnd!(gnd!), .vdd!(vdd!), .A(extDone), .B(CTRL_IDEC2_cu_custom_inst), .C(CTRL_IDEC2_cu_lui_inst), .D(CTRL_IDEC2_cu_system_inst), .Q(_2492_) );
NA3I1X1 NA3I1X1_107 ( .gnd!(gnd!), .vdd!(vdd!), .AN(_685__3_), .B(_2358_), .C(_2360_), .Q(_2493_) );
ON31X1 ON31X1_84 ( .gnd!(gnd!), .vdd!(vdd!), .A(_685__0_), .B(_685__1_), .C(_2493_), .D(_2329__bF_buf2), .Q(_2494_) );
AN31X1 AN31X1_76 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2490_), .B(_2491_), .C(_2492_), .D(_2494_), .Q(_688_) );
NO3X1 NO3X1_12 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_IDEC0_cu_alu_i_inst), .B(CTRL_IDEC0_cu_alu_r_inst), .C(CTRL_IDEC0_cu_br_inst), .Q(_2495_) );
NO2X1 NO2X1_295 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_IDEC0_cu_store_inst), .B(CTRL_IDEC0_cu_load_inst), .Q(_2496_) );
NO3X1 NO3X1_13 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_IDEC0_cu_custom_inst), .B(CTRL_IDEC0_cu_jalr_inst), .C(CTRL_IDEC0_cu_system_inst), .Q(_2497_) );
AN31X1 AN31X1_77 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2496_), .B(_2495_), .C(_2497_), .D(_2329__bF_buf3), .Q(CTRL_cu_r1_ld) );
AN21X1 AN21X1_152 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2353_), .B(_2391_), .C(_686__0_), .Q(_2498_) );
EN2X1 EN2X1_15 ( .gnd!(gnd!), .vdd!(vdd!), .A(_686__3_), .B(CTRL_IDEC1_IR_10_), .Q(_2499_) );
EN2X1 EN2X1_16 ( .gnd!(gnd!), .vdd!(vdd!), .A(_686__4_), .B(CTRL_IDEC1_IR_11_), .Q(_2500_) );
EN2X1 EN2X1_17 ( .gnd!(gnd!), .vdd!(vdd!), .A(_686__1_), .B(CTRL_IDEC1_IR_8_), .Q(_2501_) );
NA3X1 NA3X1_13 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2499_), .B(_2500_), .C(_2501_), .Q(_2502_) );
NO2X1 NO2X1_296 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_IDEC1_cu_alu_i_inst), .B(CTRL_IDEC1_cu_alu_r_inst), .Q(_2503_) );
NO3X1 NO3X1_14 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_IDEC1_cu_custom_inst_bF_buf5), .B(CTRL_IDEC1_cu_system_inst_bF_buf0), .C(CTRL_IDEC1_cu_load_inst_bF_buf2), .Q(_2504_) );
NO2X1 NO2X1_297 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_IDEC1_cu_auipc_inst_bF_buf3), .B(CTRL_IDEC1_cu_lui_inst), .Q(_2505_) );
NA3X1 NA3X1_14 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2503_), .B(_2505_), .C(_2504_), .Q(_2506_) );
AN22X1 AN22X1_70 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2391_), .B(_686__0_), .C(_686__2_), .D(_2359_), .Q(_2507_) );
ON211X1 ON211X1_108 ( .gnd!(gnd!), .vdd!(vdd!), .A(_686__2_), .B(_2359_), .C(_2507_), .D(_2506_), .Q(_2508_) );
NO3X1 NO3X1_15 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2508_), .B(_2498_), .C(_2502_), .Q(CTRL_cu_r1_src) );
NO2X1 NO2X1_298 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_IDEC0_cu_store_inst), .B(CTRL_IDEC0_cu_custom_inst), .Q(_2509_) );
AN21X1 AN21X1_153 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2495_), .B(_2509_), .C(_2329__bF_buf3), .Q(CTRL_cu_r2_ld) );
EN2X1 EN2X1_18 ( .gnd!(gnd!), .vdd!(vdd!), .A(_687__0_), .B(CTRL_IDEC1_IR_7_), .Q(_2510_) );
EN2X1 EN2X1_19 ( .gnd!(gnd!), .vdd!(vdd!), .A(_687__1_), .B(CTRL_IDEC1_IR_8_), .Q(_2511_) );
EN2X1 EN2X1_20 ( .gnd!(gnd!), .vdd!(vdd!), .A(_687__2_), .B(CTRL_IDEC1_IR_9_), .Q(_2512_) );
EN2X1 EN2X1_21 ( .gnd!(gnd!), .vdd!(vdd!), .A(_687__4_), .B(CTRL_IDEC1_IR_11_), .Q(_2513_) );
EN2X1 EN2X1_22 ( .gnd!(gnd!), .vdd!(vdd!), .A(_687__3_), .B(CTRL_IDEC1_IR_10_), .Q(_2514_) );
AND3X4 AND3X4_14 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2506_), .B(_2513_), .C(_2514_), .Q(_2515_) );
NA3I1X1 NA3I1X1_108 ( .gnd!(gnd!), .vdd!(vdd!), .AN(_687__4_), .B(_2347_), .C(_2350_), .Q(_2516_) );
AND5X2 AND5X2_1 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2510_), .B(_2511_), .C(_2512_), .D(_2516_), .E(_2515_), .Q(CTRL_cu_r2_src) );
NO2X1 NO2X1_299 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_IDEC1_cu_alu_i_inst), .B(CTRL_IDEC1_cu_jalr_inst_bF_buf4), .Q(_2517_) );
NO2X1 NO2X1_300 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_IDEC1_cu_store_inst), .B(CTRL_IDEC1_cu_load_inst_bF_buf1), .Q(_2518_) );
NA3X2 NA3X2_1 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2505_), .B(_2517_), .C(_2518_), .Q(CTRL_cu_alu_b_src) );
NO2X1 NO2X1_301 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_cu_csr_rd_s1_bF_buf2), .B(ALU_shamt_1_), .Q(_2519_) );
NA3X1 NA3X1_15 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2484_), .B(_2519_), .C(_2483_), .Q(_2520_) );
NO2X3 NO2X3_2 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2520_), .B(_2481_), .Q(CNTR_ld_cycle) );
NO2X1 NO2X1_302 ( .gnd!(gnd!), .vdd!(vdd!), .A(ALU_func7_5_bF_buf3), .B(ALU_func7_6_), .Q(_2521_) );
NA3I1X1 NA3I1X1_109 ( .gnd!(gnd!), .vdd!(vdd!), .AN(ALU_shamt_3_), .B(ALU_shamt_2_), .C(_2521_), .Q(_2522_) );
NA2X1 NA2X1_701 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2482_), .B(_2519_), .Q(_2523_) );
NO3X1 NO3X1_16 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2481_), .B(_2522_), .C(_2523_), .Q(CNTR_ld_uie) );
NO2X1 NO2X1_303 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_cu_ext_hold_bF_buf6), .B(_2475_), .Q(CTRL_cu_ld_epc) );
INX2 INX2_12 ( .gnd!(gnd!), .vdd!(vdd!), .A(rst), .Q(_2458_) );
DFRQX1 DFRQX1_129 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf30), .D(_2327_), .Q(CTRL_BR_vf) );
DFRQX1 DFRQX1_130 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf30), .D(_2328_), .Q(CTRL_BR_zf) );
DFRQX1 DFRQX1_131 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf30), .D(_2325_), .Q(CTRL_BR_sf) );
DFRQX1 DFRQX1_132 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf30), .D(_2321_), .Q(CTRL_BR_cf) );
DFRQX1 DFRQX1_133 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf48), .D(_2324_), .Q(CTRL_ISRMode) );
DFRQX1 DFRQX1_134 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf44), .D(_2326_), .Q(CTRL_TMRIF) );
DFRRQX1 DFRRQX1_157 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf48), .D(CTRL_IDEC1_cu_custom_inst_bF_buf3), .Q(_683_), .RN(_2458__bF_buf2) );
DFRRQX1 DFRRQX1_158 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf16), .D(_2323__2_), .Q(CTRL_IDEC2_IR_2_), .RN(_2458__bF_buf5) );
DFRRQX1 DFRRQX1_159 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf0), .D(_2323__3_), .Q(CTRL_IDEC2_IR_3_), .RN(_2458__bF_buf1) );
DFRSQX1 DFRSQX1_4 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf24), .D(_2323__4_), .Q(CTRL_IDEC2_IR_4_), .SN(_2458__bF_buf2) );
DFRRQX1 DFRRQX1_160 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf16), .D(_2323__5_), .Q(CTRL_IDEC2_IR_5_), .RN(_2458__bF_buf5) );
DFRRQX1 DFRRQX1_161 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf20), .D(_2323__6_), .Q(CTRL_IDEC2_IR_6_), .RN(_2458__bF_buf0) );
DFRRQX1 DFRRQX1_162 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf20), .D(_2323__7_), .Q(_685__0_), .RN(_2458__bF_buf0) );
DFRRQX1 DFRRQX1_163 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf20), .D(_2323__8_), .Q(_685__1_), .RN(_2458__bF_buf0) );
DFRRQX1 DFRRQX1_164 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf20), .D(_2323__9_), .Q(_685__2_), .RN(_2458__bF_buf0) );
DFRRQX1 DFRRQX1_165 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf16), .D(_2323__10_), .Q(_685__3_), .RN(_2458__bF_buf5) );
DFRRQX1 DFRRQX1_166 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf20), .D(_2323__11_), .Q(_685__4_), .RN(_2458__bF_buf0) );
DFRRQX1 DFRRQX1_167 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf52), .D(_2322__2_), .Q(ALU_opcode_0_), .RN(_2458__bF_buf1) );
DFRRQX1 DFRRQX1_168 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf33), .D(_2322__3_), .Q(ALU_opcode_1_), .RN(_2458__bF_buf3) );
DFRSQX2 DFRSQX2_1 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf33), .D(_2322__4_), .Q(ALU_opcode_2_), .SN(_2458__bF_buf3) );
DFRRQX2 DFRRQX2_5 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf18), .D(_2322__5_), .Q(ALU_opcode_3_), .RN(_2458__bF_buf5) );
DFRRQX2 DFRRQX2_6 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf16), .D(_2322__6_), .Q(ALU_opcode_4_), .RN(_2458__bF_buf5) );
DFRRQX1 DFRRQX1_169 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf48), .D(_2322__7_), .Q(CTRL_IDEC1_IR_7_), .RN(_2458__bF_buf4) );
DFRRQX1 DFRRQX1_170 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf20), .D(_2322__8_), .Q(CTRL_IDEC1_IR_8_), .RN(_2458__bF_buf0) );
DFRRQX1 DFRRQX1_171 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf24), .D(_2322__9_), .Q(CTRL_IDEC1_IR_9_), .RN(_2458__bF_buf2) );
DFRRQX1 DFRRQX1_172 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf16), .D(_2322__10_), .Q(CTRL_IDEC1_IR_10_), .RN(_2458__bF_buf5) );
DFRRQX1 DFRRQX1_173 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf20), .D(_2322__11_), .Q(CTRL_IDEC1_IR_11_), .RN(_2458__bF_buf4) );
DFRRQX2 DFRRQX2_7 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf33), .D(_2322__12_), .Q(_682__0_), .RN(_2458__bF_buf3) );
DFRRQX2 DFRRQX2_8 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf52), .D(_2322__13_), .Q(_682__1_), .RN(_2458__bF_buf3) );
DFRRQX4 DFRRQX4_1 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf52), .D(_2322__14_), .Q(EXT_type), .RN(_2458__bF_buf1) );
DFRRQX4 DFRRQX4_2 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf39), .D(_2322__20_), .Q(CTRL_cu_csr_rd_s1), .RN(_2458__bF_buf2) );
DFRRQX1 DFRRQX1_174 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf48), .D(_2322__21_), .Q(ALU_shamt_1_), .RN(_2458__bF_buf4) );
DFRRQX1 DFRRQX1_175 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf48), .D(_2322__22_), .Q(ALU_shamt_2_), .RN(_2458__bF_buf4) );
DFRRQX1 DFRRQX1_176 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf52), .D(_2322__23_), .Q(ALU_shamt_3_), .RN(_2458__bF_buf1) );
DFRRQX1 DFRRQX1_177 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf33), .D(_2322__24_), .Q(ALU_shamt_4_), .RN(_2458__bF_buf3) );
DFRRQX1 DFRRQX1_178 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf52), .D(_2322__25_), .Q(ALU_func7_0_), .RN(_2458__bF_buf3) );
DFRRQX1 DFRRQX1_179 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf18), .D(_2322__26_), .Q(ALU_func7_1_), .RN(_2458__bF_buf1) );
DFRRQX1 DFRRQX1_180 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf16), .D(_2322__27_), .Q(CTRL_cu_csr_rd_s2), .RN(_2458__bF_buf4) );
DFRRQX1 DFRRQX1_181 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf48), .D(_2322__28_), .Q(ALU_func7_3_), .RN(_2458__bF_buf2) );
DFRRQX1 DFRRQX1_182 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf48), .D(_2322__29_), .Q(ALU_func7_4_), .RN(_2458__bF_buf4) );
DFRRQX2 DFRRQX2_9 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf52), .D(_2322__30_), .Q(ALU_func7_5_), .RN(_2458__bF_buf1) );
DFRRQX1 DFRRQX1_183 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf48), .D(_2322__31_), .Q(ALU_func7_6_), .RN(_2458__bF_buf2) );
DFRRQX4 DFRRQX4_3 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf16), .D(_2329__bF_buf2), .Q(CTRL_cyc), .RN(_2458__bF_buf5) );
NO2X1 NO2X1_304 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_BR_vf), .B(CTRL_BR_sf), .Q(_2537_) );
AND2X2 AND2X2_70 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_BR_vf), .B(CTRL_BR_sf), .Q(_2524_) );
NO2X1 NO2X1_305 ( .gnd!(gnd!), .vdd!(vdd!), .A(_682__0_bF_buf0), .B(_682__1_bF_buf1), .Q(_2525_) );
AN211X1 AN211X1_14 ( .gnd!(gnd!), .vdd!(vdd!), .A(EXT_type_bF_buf3), .B(_2525_), .C(_2537_), .D(_2524_), .Q(_2526_) );
OR2X2 OR2X2_18 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_BR_vf), .B(CTRL_BR_sf), .Q(_2527_) );
NA2X1 NA2X1_702 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_BR_vf), .B(CTRL_BR_sf), .Q(_2528_) );
NO2I1X1 NO2I1X1_43 ( .gnd!(gnd!), .vdd!(vdd!), .AN(_682__0_bF_buf1), .B(_682__1_bF_buf4), .Q(_2529_) );
AN22X1 AN22X1_71 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2527_), .B(_2528_), .C(EXT_type_bF_buf3), .D(_2529_), .Q(_2530_) );
AND2X2 AND2X2_71 ( .gnd!(gnd!), .vdd!(vdd!), .A(_682__0_bF_buf1), .B(CTRL_BR_cf), .Q(_2531_) );
NO2X1 NO2X1_306 ( .gnd!(gnd!), .vdd!(vdd!), .A(_682__0_bF_buf1), .B(CTRL_BR_cf), .Q(_2532_) );
ON211X1 ON211X1_109 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2531_), .B(_2532_), .C(_682__1_bF_buf1), .D(EXT_type_bF_buf3), .Q(_2533_) );
INX1 INX1_188 ( .gnd!(gnd!), .vdd!(vdd!), .A(EXT_type_bF_buf5), .Q(_2534_) );
ON21X1 ON21X1_303 ( .gnd!(gnd!), .vdd!(vdd!), .A(_682__0_bF_buf1), .B(_682__1_bF_buf1), .C(CTRL_BR_zf), .Q(_2535_) );
ON211X1 ON211X1_110 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2529_), .B(CTRL_BR_zf), .C(_2534_), .D(_2535_), .Q(_2536_) );
ON211X1 ON211X1_111 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2526_), .B(_2530_), .C(_2536_), .D(_2533_), .Q(CTRL_BR_taken) );
NA2I1X1 NA2I1X1_100 ( .gnd!(gnd!), .vdd!(vdd!), .AN(CTRL_IDEC0_IR_4_), .B(CTRL_IDEC0_IR_5_), .Q(_2538_) );
NO2X1 NO2X1_307 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_IDEC0_IR_2_), .B(CTRL_IDEC0_IR_3_), .Q(_2539_) );
NA2X1 NA2X1_703 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2539_), .B(CTRL_IDEC0_IR_6_), .Q(_2540_) );
NO2X1 NO2X1_308 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2538_), .B(_2540_), .Q(CTRL_IDEC0_cu_br_inst) );
NA3I1X1 NA3I1X1_110 ( .gnd!(gnd!), .vdd!(vdd!), .AN(CTRL_IDEC0_IR_3_), .B(CTRL_IDEC0_IR_2_), .C(CTRL_IDEC0_IR_6_), .Q(_2541_) );
NO2X1 NO2X1_309 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2538_), .B(_2541_), .Q(CTRL_IDEC0_cu_jalr_inst) );
NA2I1X1 NA2I1X1_101 ( .gnd!(gnd!), .vdd!(vdd!), .AN(CTRL_IDEC0_IR_6_), .B(_2539_), .Q(_2542_) );
NA2I1X1 NA2I1X1_102 ( .gnd!(gnd!), .vdd!(vdd!), .AN(CTRL_IDEC0_IR_5_), .B(CTRL_IDEC0_IR_4_), .Q(_2543_) );
NO2X1 NO2X1_310 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2543_), .B(_2542_), .Q(CTRL_IDEC0_cu_alu_i_inst) );
NA2X1 NA2X1_704 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_IDEC0_IR_5_), .B(CTRL_IDEC0_IR_4_), .Q(_2544_) );
NO2X1 NO2X1_311 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2544_), .B(_2542_), .Q(CTRL_IDEC0_cu_alu_r_inst) );
OR2X2 OR2X2_19 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_IDEC0_IR_5_), .B(CTRL_IDEC0_IR_4_), .Q(_2545_) );
NO2X1 NO2X1_312 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2545_), .B(_2542_), .Q(CTRL_IDEC0_cu_load_inst) );
NO2X1 NO2X1_313 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2538_), .B(_2542_), .Q(CTRL_IDEC0_cu_store_inst) );
NO2X1 NO2X1_314 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2545_), .B(_2541_), .Q(CTRL_IDEC0_cu_custom_inst) );
NO2X1 NO2X1_315 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2544_), .B(_2540_), .Q(CTRL_IDEC0_cu_system_inst) );
NA2I1X1 NA2I1X1_103 ( .gnd!(gnd!), .vdd!(vdd!), .AN(ALU_opcode_2_), .B(ALU_opcode_3_), .Q(_2546_) );
NO2X1 NO2X1_316 ( .gnd!(gnd!), .vdd!(vdd!), .A(ALU_opcode_0_), .B(ALU_opcode_1_), .Q(_2547_) );
NA2X1 NA2X1_705 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2547_), .B(ALU_opcode_4_), .Q(_2548_) );
NO2X1 NO2X1_317 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2546_), .B(_2548_), .Q(CTRL_IDEC1_cu_br_inst) );
NA3I1X1 NA3I1X1_111 ( .gnd!(gnd!), .vdd!(vdd!), .AN(ALU_opcode_2_), .B(ALU_opcode_3_), .C(ALU_opcode_4_), .Q(_2549_) );
NA2X1 NA2X1_706 ( .gnd!(gnd!), .vdd!(vdd!), .A(ALU_opcode_0_), .B(ALU_opcode_1_), .Q(_2550_) );
NO2X1 NO2X1_318 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2550_), .B(_2549_), .Q(CTRL_IDEC1_cu_jal_inst) );
NA3I1X1 NA3I1X1_112 ( .gnd!(gnd!), .vdd!(vdd!), .AN(ALU_opcode_1_), .B(ALU_opcode_0_), .C(ALU_opcode_4_), .Q(_2551_) );
NO2X2 NO2X2_4 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2546_), .B(_2551_), .Q(CTRL_IDEC1_cu_jalr_inst) );
NA2I1X1 NA2I1X1_104 ( .gnd!(gnd!), .vdd!(vdd!), .AN(ALU_opcode_4_), .B(_2547_), .Q(_2552_) );
NA2I1X1 NA2I1X1_105 ( .gnd!(gnd!), .vdd!(vdd!), .AN(ALU_opcode_3_), .B(ALU_opcode_2_), .Q(_2553_) );
NO2X1 NO2X1_319 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2553_), .B(_2552_), .Q(CTRL_IDEC1_cu_alu_i_inst) );
NA2X1 NA2X1_707 ( .gnd!(gnd!), .vdd!(vdd!), .A(ALU_opcode_3_), .B(ALU_opcode_2_), .Q(_2554_) );
NO2X1 NO2X1_320 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2554_), .B(_2552_), .Q(CTRL_IDEC1_cu_alu_r_inst) );
OR2X2 OR2X2_20 ( .gnd!(gnd!), .vdd!(vdd!), .A(ALU_opcode_3_), .B(ALU_opcode_2_), .Q(_2555_) );
NO2X2 NO2X2_5 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2555_), .B(_2552_), .Q(CTRL_IDEC1_cu_load_inst) );
NO2X1 NO2X1_321 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2546_), .B(_2552_), .Q(CTRL_IDEC1_cu_store_inst) );
NA3I2X1 NA3I2X1_26 ( .gnd!(gnd!), .vdd!(vdd!), .AN(ALU_opcode_1_), .BN(ALU_opcode_4_), .C(ALU_opcode_0_), .Q(_2556_) );
NO2X1 NO2X1_322 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2554_), .B(_2556_), .Q(CTRL_IDEC1_cu_lui_inst) );
NO2X2 NO2X2_6 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2553_), .B(_2556_), .Q(CTRL_IDEC1_cu_auipc_inst) );
NO2X2 NO2X2_7 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2555_), .B(_2551_), .Q(CTRL_IDEC1_cu_custom_inst) );
NO2X3 NO2X3_3 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2554_), .B(_2548_), .Q(CTRL_IDEC1_cu_system_inst) );
NA2I1X1 NA2I1X1_106 ( .gnd!(gnd!), .vdd!(vdd!), .AN(CTRL_IDEC2_IR_4_), .B(CTRL_IDEC2_IR_5_), .Q(_2557_) );
NO2X1 NO2X1_323 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_IDEC2_IR_2_), .B(CTRL_IDEC2_IR_3_), .Q(_2558_) );
NA2X1 NA2X1_708 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2558_), .B(CTRL_IDEC2_IR_6_), .Q(_2559_) );
NA3I1X1 NA3I1X1_113 ( .gnd!(gnd!), .vdd!(vdd!), .AN(CTRL_IDEC2_IR_4_), .B(CTRL_IDEC2_IR_5_), .C(CTRL_IDEC2_IR_6_), .Q(_2560_) );
NA2X1 NA2X1_709 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_IDEC2_IR_2_), .B(CTRL_IDEC2_IR_3_), .Q(_2561_) );
NO2X1 NO2X1_324 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2561_), .B(_2560_), .Q(CTRL_IDEC2_cu_jal_inst) );
NA3I1X1 NA3I1X1_114 ( .gnd!(gnd!), .vdd!(vdd!), .AN(CTRL_IDEC2_IR_3_), .B(CTRL_IDEC2_IR_2_), .C(CTRL_IDEC2_IR_6_), .Q(_2562_) );
NO2X1 NO2X1_325 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2557_), .B(_2562_), .Q(CTRL_IDEC2_cu_jalr_inst) );
NA2I1X1 NA2I1X1_107 ( .gnd!(gnd!), .vdd!(vdd!), .AN(CTRL_IDEC2_IR_6_), .B(_2558_), .Q(_2563_) );
NA2I1X1 NA2I1X1_108 ( .gnd!(gnd!), .vdd!(vdd!), .AN(CTRL_IDEC2_IR_5_), .B(CTRL_IDEC2_IR_4_), .Q(_2564_) );
NO2X1 NO2X1_326 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2564_), .B(_2563_), .Q(CTRL_IDEC2_cu_alu_i_inst) );
NA2X1 NA2X1_710 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_IDEC2_IR_5_), .B(CTRL_IDEC2_IR_4_), .Q(_2565_) );
NO2X1 NO2X1_327 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2565_), .B(_2563_), .Q(CTRL_IDEC2_cu_alu_r_inst) );
OR2X2 OR2X2_21 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_IDEC2_IR_5_), .B(CTRL_IDEC2_IR_4_), .Q(_2566_) );
NO2X1 NO2X1_328 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2566_), .B(_2563_), .Q(CTRL_IDEC2_cu_load_inst) );
NA3I2X1 NA3I2X1_27 ( .gnd!(gnd!), .vdd!(vdd!), .AN(CTRL_IDEC2_IR_3_), .BN(CTRL_IDEC2_IR_6_), .C(CTRL_IDEC2_IR_2_), .Q(_2567_) );
NO2X1 NO2X1_329 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2565_), .B(_2567_), .Q(CTRL_IDEC2_cu_lui_inst) );
NO2X1 NO2X1_330 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2564_), .B(_2567_), .Q(CTRL_IDEC2_cu_auipc_inst) );
NO2X1 NO2X1_331 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2566_), .B(_2562_), .Q(CTRL_IDEC2_cu_custom_inst) );
NO2X1 NO2X1_332 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2565_), .B(_2559_), .Q(CTRL_IDEC2_cu_system_inst) );
INX1 INX1_189 ( .gnd!(gnd!), .vdd!(vdd!), .A(bdo[8]), .Q(_2571_) );
NO2X1 NO2X1_333 ( .gnd!(gnd!), .vdd!(vdd!), .A(_682__1_bF_buf4), .B(_682__0_bF_buf2), .Q(_2572_) );
NA2X1 NA2X1_711 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2572_), .B(bdo[7]), .Q(_2573_) );
ON22X1 ON22X1_76 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2573_), .B(EXT_type_bF_buf5), .C(_2571_), .D(_2572_), .Q(EXT_do_8_) );
INX1 INX1_190 ( .gnd!(gnd!), .vdd!(vdd!), .A(bdo[9]), .Q(_2574_) );
ON22X1 ON22X1_77 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2573_), .B(EXT_type_bF_buf5), .C(_2574_), .D(_2572_), .Q(EXT_do_9_) );
INX1 INX1_191 ( .gnd!(gnd!), .vdd!(vdd!), .A(bdo[10]), .Q(_2575_) );
ON22X1 ON22X1_78 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2573_), .B(EXT_type_bF_buf0), .C(_2575_), .D(_2572_), .Q(EXT_do_10_) );
INX1 INX1_192 ( .gnd!(gnd!), .vdd!(vdd!), .A(bdo[11]), .Q(_2576_) );
ON22X1 ON22X1_79 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2573_), .B(EXT_type_bF_buf5), .C(_2576_), .D(_2572_), .Q(EXT_do_11_) );
INX1 INX1_193 ( .gnd!(gnd!), .vdd!(vdd!), .A(bdo[12]), .Q(_2577_) );
ON22X1 ON22X1_80 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2573_), .B(EXT_type_bF_buf5), .C(_2577_), .D(_2572_), .Q(EXT_do_12_) );
INX1 INX1_194 ( .gnd!(gnd!), .vdd!(vdd!), .A(bdo[13]), .Q(_2578_) );
ON22X1 ON22X1_81 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2573_), .B(EXT_type_bF_buf5), .C(_2578_), .D(_2572_), .Q(EXT_do_13_) );
INX1 INX1_195 ( .gnd!(gnd!), .vdd!(vdd!), .A(bdo[14]), .Q(_2579_) );
ON22X1 ON22X1_82 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2573_), .B(EXT_type_bF_buf5), .C(_2579_), .D(_2572_), .Q(EXT_do_14_) );
INX1 INX1_196 ( .gnd!(gnd!), .vdd!(vdd!), .A(bdo[15]), .Q(_2580_) );
ON22X1 ON22X1_83 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2573_), .B(EXT_type_bF_buf0), .C(_2580_), .D(_2572_), .Q(EXT_do_15_) );
OR2X2 OR2X2_22 ( .gnd!(gnd!), .vdd!(vdd!), .A(_682__1_bF_buf0), .B(_682__0_bF_buf2), .Q(_2581_) );
NA2I1X2 NA2I1X2_2 ( .gnd!(gnd!), .vdd!(vdd!), .AN(EXT_type_bF_buf0), .B(bdo[7]), .Q(_2582_) );
NA2I1X1 NA2I1X1_109 ( .gnd!(gnd!), .vdd!(vdd!), .AN(_682__1_bF_buf0), .B(_682__0_bF_buf2), .Q(_2583_) );
NA2X1 NA2X1_712 ( .gnd!(gnd!), .vdd!(vdd!), .A(_682__1_bF_buf2), .B(bdo[16]), .Q(_2584_) );
NA2I1X2 NA2I1X2_3 ( .gnd!(gnd!), .vdd!(vdd!), .AN(EXT_type_bF_buf0), .B(bdo[15]), .Q(_2585_) );
ON221X1 ON221X1_5 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2583_), .B(_2585_), .C(_2582_), .D(_2581_), .E(_2584_), .Q(EXT_do_16_) );
NA2X1 NA2X1_713 ( .gnd!(gnd!), .vdd!(vdd!), .A(_682__1_bF_buf0), .B(bdo[17]), .Q(_2586_) );
ON221X1 ON221X1_6 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2583_), .B(_2585_), .C(_2582_), .D(_2581_), .E(_2586_), .Q(EXT_do_17_) );
NA2X1 NA2X1_714 ( .gnd!(gnd!), .vdd!(vdd!), .A(_682__1_bF_buf0), .B(bdo[18]), .Q(_2587_) );
ON221X1 ON221X1_7 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2583_), .B(_2585_), .C(_2582_), .D(_2581_), .E(_2587_), .Q(EXT_do_18_) );
NA2X1 NA2X1_715 ( .gnd!(gnd!), .vdd!(vdd!), .A(_682__1_bF_buf3), .B(bdo[19]), .Q(_2588_) );
ON221X1 ON221X1_8 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2583_), .B(_2585_), .C(_2582_), .D(_2581_), .E(_2588_), .Q(EXT_do_19_) );
NA2X1 NA2X1_716 ( .gnd!(gnd!), .vdd!(vdd!), .A(_682__1_bF_buf3), .B(bdo[20]), .Q(_2589_) );
ON221X1 ON221X1_9 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2583_), .B(_2585_), .C(_2582_), .D(_2581_), .E(_2589_), .Q(EXT_do_20_) );
NA2X1 NA2X1_717 ( .gnd!(gnd!), .vdd!(vdd!), .A(_682__1_bF_buf2), .B(bdo[21]), .Q(_2590_) );
ON221X1 ON221X1_10 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2583_), .B(_2585_), .C(_2582_), .D(_2581_), .E(_2590_), .Q(EXT_do_21_) );
NA2X1 NA2X1_718 ( .gnd!(gnd!), .vdd!(vdd!), .A(_682__1_bF_buf2), .B(bdo[22]), .Q(_2591_) );
ON221X1 ON221X1_11 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2583_), .B(_2585_), .C(_2582_), .D(_2581_), .E(_2591_), .Q(EXT_do_22_) );
NA2X1 NA2X1_719 ( .gnd!(gnd!), .vdd!(vdd!), .A(_682__1_bF_buf2), .B(bdo[23]), .Q(_2592_) );
ON221X1 ON221X1_12 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2583_), .B(_2585_), .C(_2582_), .D(_2581_), .E(_2592_), .Q(EXT_do_23_) );
NA2X1 NA2X1_720 ( .gnd!(gnd!), .vdd!(vdd!), .A(_682__1_bF_buf3), .B(bdo[24]), .Q(_2593_) );
ON221X1 ON221X1_13 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2583_), .B(_2585_), .C(_2582_), .D(_2581_), .E(_2593_), .Q(EXT_do_24_) );
NA2X1 NA2X1_721 ( .gnd!(gnd!), .vdd!(vdd!), .A(_682__1_bF_buf3), .B(bdo[25]), .Q(_2594_) );
ON221X1 ON221X1_14 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2583_), .B(_2585_), .C(_2582_), .D(_2581_), .E(_2594_), .Q(EXT_do_25_) );
NA2X1 NA2X1_722 ( .gnd!(gnd!), .vdd!(vdd!), .A(_682__1_bF_buf4), .B(bdo[26]), .Q(_2595_) );
ON221X1 ON221X1_15 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2583_), .B(_2585_), .C(_2582_), .D(_2581_), .E(_2595_), .Q(EXT_do_26_) );
NA2X1 NA2X1_723 ( .gnd!(gnd!), .vdd!(vdd!), .A(_682__1_bF_buf3), .B(bdo[27]), .Q(_2596_) );
ON221X1 ON221X1_16 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2583_), .B(_2585_), .C(_2582_), .D(_2581_), .E(_2596_), .Q(EXT_do_27_) );
NA2X1 NA2X1_724 ( .gnd!(gnd!), .vdd!(vdd!), .A(_682__1_bF_buf0), .B(bdo[28]), .Q(_2597_) );
ON221X1 ON221X1_17 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2583_), .B(_2585_), .C(_2582_), .D(_2581_), .E(_2597_), .Q(EXT_do_28_) );
NA2X1 NA2X1_725 ( .gnd!(gnd!), .vdd!(vdd!), .A(_682__1_bF_buf3), .B(bdo[29]), .Q(_2568_) );
ON221X1 ON221X1_18 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2583_), .B(_2585_), .C(_2582_), .D(_2581_), .E(_2568_), .Q(EXT_do_29_) );
NA2X1 NA2X1_726 ( .gnd!(gnd!), .vdd!(vdd!), .A(_682__1_bF_buf0), .B(bdo[30]), .Q(_2569_) );
ON221X1 ON221X1_19 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2583_), .B(_2585_), .C(_2582_), .D(_2581_), .E(_2569_), .Q(EXT_do_30_) );
NA2X1 NA2X1_727 ( .gnd!(gnd!), .vdd!(vdd!), .A(_682__1_bF_buf3), .B(bdo[31]), .Q(_2570_) );
ON221X1 ON221X1_20 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2583_), .B(_2585_), .C(_2582_), .D(_2581_), .E(_2570_), .Q(EXT_do_31_) );
INX1 INX1_197 ( .gnd!(gnd!), .vdd!(vdd!), .A(_687__0_), .Q(_2614_) );
NA2X1 NA2X1_728 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_IDEC0_IR_2_), .B(CTRL_IDEC0_IR_4_), .Q(_2615_) );
NO3X1 NO3X1_17 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2615_), .B(CTRL_IDEC0_IR_3_), .C(CTRL_IDEC0_IR_6_), .Q(_2616_) );
NO2X1 NO2X1_334 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_IDEC0_IR_2_), .B(CTRL_IDEC0_IR_3_), .Q(_2617_) );
NA3I1X1 NA3I1X1_115 ( .gnd!(gnd!), .vdd!(vdd!), .AN(CTRL_IDEC0_IR_4_), .B(CTRL_IDEC0_IR_5_), .C(_2617_), .Q(_2618_) );
NA2I1X1 NA2I1X1_110 ( .gnd!(gnd!), .vdd!(vdd!), .AN(CTRL_IDEC0_IR_4_), .B(CTRL_IDEC0_IR_5_), .Q(_2619_) );
NA3X1 NA3X1_16 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_IDEC0_IR_2_), .B(CTRL_IDEC0_IR_3_), .C(CTRL_IDEC0_IR_6_), .Q(_2620_) );
ON21X1 ON21X1_304 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2619_), .B(_2620_), .C(_2618_), .Q(_2621_) );
NA2I1X1 NA2I1X1_111 ( .gnd!(gnd!), .vdd!(vdd!), .AN(CTRL_IDEC0_IR_6_), .B(CTRL_IDEC0_IR_7_), .Q(_2622_) );
ON32X1 ON32X1_5 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2614_), .B(_2616_), .C(_2621_), .D(_2618_), .E(_2622_), .Q(IMM_0_) );
INX1 INX1_198 ( .gnd!(gnd!), .vdd!(vdd!), .A(_687__1_), .Q(_2623_) );
NO3X1 NO3X1_18 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2619_), .B(CTRL_IDEC0_IR_2_), .C(CTRL_IDEC0_IR_3_), .Q(_2624_) );
NA2X1 NA2X1_729 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2624_), .B(CTRL_IDEC0_IR_8_), .Q(_2625_) );
NO2X1 NO2X1_335 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_IDEC0_IR_3_), .B(CTRL_IDEC0_IR_6_), .Q(_2626_) );
NA2I1X1 NA2I1X1_112 ( .gnd!(gnd!), .vdd!(vdd!), .AN(_2615_), .B(_2626_), .Q(_2627_) );
NO2X1 NO2X1_336 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2620_), .B(_2619_), .Q(_2628_) );
AN21X1 AN21X1_154 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2627_), .B(_2618_), .C(_2628_), .Q(_2629_) );
ON21X1 ON21X1_305 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2629_), .B(_2623_), .C(_2625_), .Q(IMM_1_) );
INX1 INX1_199 ( .gnd!(gnd!), .vdd!(vdd!), .A(_687__2_), .Q(_2630_) );
NA2X1 NA2X1_730 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2624_), .B(CTRL_IDEC0_IR_9_), .Q(_2631_) );
ON21X1 ON21X1_306 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2629_), .B(_2630_), .C(_2631_), .Q(IMM_2_) );
INX1 INX1_200 ( .gnd!(gnd!), .vdd!(vdd!), .A(_687__3_), .Q(_2632_) );
NA2X1 NA2X1_731 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2624_), .B(CTRL_IDEC0_IR_10_), .Q(_2633_) );
ON21X1 ON21X1_307 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2629_), .B(_2632_), .C(_2633_), .Q(IMM_3_) );
INX1 INX1_201 ( .gnd!(gnd!), .vdd!(vdd!), .A(_687__4_), .Q(_2634_) );
NA2X1 NA2X1_732 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2624_), .B(CTRL_IDEC0_IR_11_), .Q(_2635_) );
ON21X1 ON21X1_308 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2629_), .B(_2634_), .C(_2635_), .Q(IMM_4_) );
AND2X2 AND2X2_72 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2627_), .B(CTRL_IDEC0_IR_25_), .Q(IMM_5_) );
AND2X2 AND2X2_73 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2627_), .B(CTRL_IDEC0_IR_26_), .Q(IMM_6_) );
AND2X2 AND2X2_74 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2627_), .B(CTRL_IDEC0_IR_27_), .Q(IMM_7_) );
AND2X2 AND2X2_75 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2627_), .B(CTRL_IDEC0_IR_28_), .Q(IMM_8_) );
AND2X2 AND2X2_76 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2627_), .B(CTRL_IDEC0_IR_29_), .Q(IMM_9_) );
AND2X2 AND2X2_77 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2627_), .B(CTRL_IDEC0_IR_30_), .Q(IMM_10_) );
INX1 INX1_202 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_IDEC0_IR_31_), .Q(_2636_) );
ON32X1 ON32X1_6 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_IDEC0_IR_3_), .B(CTRL_IDEC0_IR_6_), .C(_2615_), .D(_2620_), .E(_2619_), .Q(_2637_) );
NA2X1 NA2X1_733 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2628_), .B(_687__0_), .Q(_2638_) );
MU2X1 MU2X1_218 ( .gnd!(gnd!), .vdd!(vdd!), .IN0(CTRL_IDEC0_IR_31_), .IN1(CTRL_IDEC0_IR_7_), .Q(_2639_), .S(CTRL_IDEC0_IR_6_) );
NA2X1 NA2X1_734 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2624_), .B(_2639_), .Q(_2640_) );
ON311X1 ON311X1_8 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2636_), .B(_2624_), .C(_2637_), .D(_2638_), .E(_2640_), .Q(IMM_11_) );
NA2X1 NA2X1_735 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2637_), .B(CTRL_IDEC0_IR_12_), .Q(_2598_) );
NA3I1X1 NA3I1X1_116 ( .gnd!(gnd!), .vdd!(vdd!), .AN(_2619_), .B(CTRL_IDEC0_IR_31_), .C(_2617_), .Q(_2599_) );
ON311X1 ON311X1_9 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2636_), .B(_2616_), .C(_2621_), .D(_2599_), .E(_2598_), .Q(IMM_12_) );
NA2X1 NA2X1_736 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2637_), .B(CTRL_IDEC0_IR_13_), .Q(_2600_) );
ON311X1 ON311X1_10 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2636_), .B(_2616_), .C(_2621_), .D(_2599_), .E(_2600_), .Q(IMM_13_) );
NA2X1 NA2X1_737 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2637_), .B(CTRL_IDEC0_IR_14_), .Q(_2601_) );
ON311X1 ON311X1_11 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2636_), .B(_2616_), .C(_2621_), .D(_2599_), .E(_2601_), .Q(IMM_14_) );
NA2X1 NA2X1_738 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2637_), .B(_686__0_), .Q(_2602_) );
ON311X1 ON311X1_12 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2636_), .B(_2616_), .C(_2621_), .D(_2599_), .E(_2602_), .Q(IMM_15_) );
NA2X1 NA2X1_739 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2637_), .B(_686__1_), .Q(_2603_) );
ON311X1 ON311X1_13 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2636_), .B(_2616_), .C(_2621_), .D(_2599_), .E(_2603_), .Q(IMM_16_) );
NA2X1 NA2X1_740 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2637_), .B(_686__2_), .Q(_2604_) );
ON311X1 ON311X1_14 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2636_), .B(_2616_), .C(_2621_), .D(_2599_), .E(_2604_), .Q(IMM_17_) );
NA2X1 NA2X1_741 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2637_), .B(_686__3_), .Q(_2605_) );
ON311X1 ON311X1_15 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2636_), .B(_2616_), .C(_2621_), .D(_2599_), .E(_2605_), .Q(IMM_18_) );
NA2X1 NA2X1_742 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2637_), .B(_686__4_), .Q(_2606_) );
ON311X1 ON311X1_16 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2636_), .B(_2616_), .C(_2621_), .D(_2599_), .E(_2606_), .Q(IMM_19_) );
NA2X1 NA2X1_743 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2627_), .B(CTRL_IDEC0_IR_31_), .Q(_2607_) );
ON21X1 ON21X1_309 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2614_), .B(_2627_), .C(_2607_), .Q(IMM_20_) );
ON21X1 ON21X1_310 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2623_), .B(_2627_), .C(_2607_), .Q(IMM_21_) );
ON21X1 ON21X1_311 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2630_), .B(_2627_), .C(_2607_), .Q(IMM_22_) );
ON21X1 ON21X1_312 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2632_), .B(_2627_), .C(_2607_), .Q(IMM_23_) );
ON21X1 ON21X1_313 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2634_), .B(_2627_), .C(_2607_), .Q(IMM_24_) );
NA2X1 NA2X1_744 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2616_), .B(CTRL_IDEC0_IR_25_), .Q(_2608_) );
NA2X1 NA2X1_745 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2607_), .B(_2608_), .Q(IMM_25_) );
NA2X1 NA2X1_746 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2616_), .B(CTRL_IDEC0_IR_26_), .Q(_2609_) );
NA2X1 NA2X1_747 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2607_), .B(_2609_), .Q(IMM_26_) );
NA2X1 NA2X1_748 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2616_), .B(CTRL_IDEC0_IR_27_), .Q(_2610_) );
NA2X1 NA2X1_749 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2607_), .B(_2610_), .Q(IMM_27_) );
NA2X1 NA2X1_750 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2616_), .B(CTRL_IDEC0_IR_28_), .Q(_2611_) );
NA2X1 NA2X1_751 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2607_), .B(_2611_), .Q(IMM_28_) );
NA2X1 NA2X1_752 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2616_), .B(CTRL_IDEC0_IR_29_), .Q(_2612_) );
NA2X1 NA2X1_753 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2607_), .B(_2612_), .Q(IMM_29_) );
NA2X1 NA2X1_754 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2616_), .B(CTRL_IDEC0_IR_30_), .Q(_2613_) );
NA2X1 NA2X1_755 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2607_), .B(_2613_), .Q(IMM_30_) );
INX2 INX2_13 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_cu_ld_epc), .Q(_2643_) );
INX1 INX1_203 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_cu_pc_s2_bF_buf2), .Q(_2644_) );
NO2X1 NO2X1_337 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_IDEC1_cu_jalr_inst_bF_buf3), .B(CTRL_cu_sel_epc), .Q(_2645_) );
NA2X1 NA2X1_756 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2644_), .B(_2645_), .Q(_2646_) );
INX2 INX2_14 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2646__bF_buf0), .Q(_2647_) );
NA2X1 NA2X1_757 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_cu_pc_s2_bF_buf2), .B(I1_0_), .Q(_2648_) );
ON21X1 ON21X1_314 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_cu_pc_s2_bF_buf1), .B(CTRL_cu_pc_s3_bF_buf1), .C(PC1_0_), .Q(_2649_) );
NO2X4 NO2X4_1 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_cu_pc_s2_bF_buf4), .B(CTRL_cu_pc_s3_bF_buf2), .Q(_2650_) );
NA2X1 NA2X1_758 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2650__bF_buf6), .B(PC_0_), .Q(_2651_) );
AN21X1 AN21X1_155 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2651_), .B(_2649_), .C(_2648_), .Q(_2652_) );
AND2X2 AND2X2_78 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_cu_pc_s2_bF_buf1), .B(I1_0_), .Q(_2653_) );
NA2X1 NA2X1_759 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2651_), .B(_2649_), .Q(_2654_) );
NO2X1 NO2X1_338 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2653_), .B(_2654_), .Q(_2655_) );
NA2X1 NA2X1_760 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_IDEC1_cu_jalr_inst_bF_buf4), .B(ALU_r_0_), .Q(_2656_) );
ON31X1 ON31X1_85 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_IDEC1_cu_jalr_inst_bF_buf5), .B(_2652_), .C(_2655_), .D(_2656_), .Q(_2657_) );
MU2X1 MU2X1_219 ( .gnd!(gnd!), .vdd!(vdd!), .IN0(_2657_), .IN1(PC_0_), .Q(_2658_), .S(_2647__bF_buf2) );
MU2X1 MU2X1_220 ( .gnd!(gnd!), .vdd!(vdd!), .IN0(_2658_), .IN1(PCU_ePC_0_), .Q(_2642__0_), .S(_2643__bF_buf5) );
NA2X1 NA2X1_761 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_cu_pc_s2_bF_buf2), .B(I1_1_), .Q(_2659_) );
ON21X1 ON21X1_315 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_cu_pc_s2_bF_buf1), .B(CTRL_cu_pc_s3_bF_buf3), .C(PC1_1_), .Q(_2660_) );
NA2X1 NA2X1_762 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2650__bF_buf6), .B(PC_1_), .Q(_2661_) );
NA3X1 NA3X1_17 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2659_), .B(_2660_), .C(_2661_), .Q(_2662_) );
AND2X2 AND2X2_79 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_cu_pc_s2_bF_buf3), .B(I1_1_), .Q(_2663_) );
NA2X1 NA2X1_763 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2661_), .B(_2660_), .Q(_2664_) );
NA2X1 NA2X1_764 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2664_), .B(_2663_), .Q(_2665_) );
NA2X1 NA2X1_765 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2665_), .B(_2662_), .Q(_2666_) );
EN2X1 EN2X1_23 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2666_), .B(_2652_), .Q(_2667_) );
MU2X1 MU2X1_221 ( .gnd!(gnd!), .vdd!(vdd!), .IN0(_2667_), .IN1(ALU_r_1_), .Q(_2668_), .S(CTRL_IDEC1_cu_jalr_inst_bF_buf3) );
MU2X1 MU2X1_222 ( .gnd!(gnd!), .vdd!(vdd!), .IN0(_2668_), .IN1(PC_1_), .Q(_2669_), .S(_2647__bF_buf1) );
MU2X1 MU2X1_223 ( .gnd!(gnd!), .vdd!(vdd!), .IN0(_2669_), .IN1(PCU_ePC_1_), .Q(_2642__1_), .S(_2643__bF_buf1) );
AN21X1 AN21X1_156 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2661_), .B(_2660_), .C(_2659_), .Q(_2670_) );
AN21X1 AN21X1_157 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2652_), .B(_2662_), .C(_2670_), .Q(_2671_) );
NA2I1X1 NA2I1X1_113 ( .gnd!(gnd!), .vdd!(vdd!), .AN(I1_2_), .B(CTRL_cu_pc_s2_bF_buf6), .Q(_2672_) );
NO3I1X1 NO3I1X1_3 ( .gnd!(gnd!), .vdd!(vdd!), .AN(PC_2_), .B(CTRL_cu_pc_s2_bF_buf1), .C(CTRL_cu_pc_s3_bF_buf3), .Q(_2673_) );
OA21X4 OA21X4_1 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_cu_pc_s2_bF_buf1), .B(CTRL_cu_pc_s3_bF_buf1), .C(PC1_2_), .Q(_2674_) );
ON21X1 ON21X1_316 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2674_), .B(_2673_), .C(_2672_), .Q(_2675_) );
NO2I1X1 NO2I1X1_44 ( .gnd!(gnd!), .vdd!(vdd!), .AN(CTRL_cu_pc_s2_bF_buf6), .B(I1_2_), .Q(_2676_) );
NA2X1 NA2X1_766 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2650__bF_buf2), .B(PC_2_), .Q(_2677_) );
ON21X1 ON21X1_317 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_cu_pc_s2_bF_buf1), .B(CTRL_cu_pc_s3_bF_buf1), .C(PC1_2_), .Q(_2678_) );
NA3X1 NA3X1_18 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2676_), .B(_2678_), .C(_2677_), .Q(_2679_) );
NA2X1 NA2X1_767 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2675_), .B(_2679_), .Q(_2680_) );
AND2X2 AND2X2_80 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2671_), .B(_2680_), .Q(_2681_) );
NO2X1 NO2X1_339 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2680_), .B(_2671_), .Q(_2682_) );
NA2X1 NA2X1_768 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_IDEC1_cu_jalr_inst_bF_buf4), .B(ALU_r_2_), .Q(_2683_) );
ON31X1 ON31X1_86 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_IDEC1_cu_jalr_inst_bF_buf5), .B(_2682_), .C(_2681_), .D(_2683_), .Q(_2684_) );
MU2X1 MU2X1_224 ( .gnd!(gnd!), .vdd!(vdd!), .IN0(_2684_), .IN1(PC_2_), .Q(_2685_), .S(_2647__bF_buf0) );
MU2X1 MU2X1_225 ( .gnd!(gnd!), .vdd!(vdd!), .IN0(_2685_), .IN1(PCU_ePC_2_), .Q(_2642__2_), .S(_2643__bF_buf1) );
INX1 INX1_204 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_IDEC1_cu_jalr_inst_bF_buf2), .Q(_2686_) );
NO2X1 NO2X1_340 ( .gnd!(gnd!), .vdd!(vdd!), .A(ALU_r_3_), .B(_2686__bF_buf3), .Q(_2687_) );
NA2X1 NA2X1_769 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_cu_pc_s2_bF_buf3), .B(I1_3_), .Q(_2688_) );
OA21X4 OA21X4_2 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_cu_pc_s2_bF_buf6), .B(CTRL_cu_pc_s3_bF_buf3), .C(PC1_3_), .Q(_2689_) );
NO3I1X1 NO3I1X1_4 ( .gnd!(gnd!), .vdd!(vdd!), .AN(PC_3_), .B(CTRL_cu_pc_s2_bF_buf6), .C(CTRL_cu_pc_s3_bF_buf1), .Q(_2690_) );
ON21X1 ON21X1_318 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2689_), .B(_2690_), .C(_2688_), .Q(_2691_) );
ON21X1 ON21X1_319 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_cu_pc_s2_bF_buf6), .B(CTRL_cu_pc_s3_bF_buf3), .C(PC1_3_), .Q(_2692_) );
NA2X1 NA2X1_770 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2650__bF_buf2), .B(PC_3_), .Q(_2693_) );
NA3I1X1 NA3I1X1_117 ( .gnd!(gnd!), .vdd!(vdd!), .AN(_2688_), .B(_2692_), .C(_2693_), .Q(_2694_) );
NA2X1 NA2X1_771 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2691_), .B(_2694_), .Q(_2695_) );
AN21X1 AN21X1_158 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2677_), .B(_2678_), .C(_2676_), .Q(_2696_) );
NO2X1 NO2X1_341 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2696_), .B(_2682_), .Q(_2697_) );
NA2X1 NA2X1_772 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2697_), .B(_2695_), .Q(_2698_) );
OR2X2 OR2X2_23 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2697_), .B(_2695_), .Q(_2699_) );
AN31X1 AN31X1_78 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2686__bF_buf3), .B(_2698_), .C(_2699_), .D(_2687_), .Q(_2700_) );
MU2X1 MU2X1_226 ( .gnd!(gnd!), .vdd!(vdd!), .IN0(_2700_), .IN1(PC_3_), .Q(_2701_), .S(_2647__bF_buf3) );
MU2X1 MU2X1_227 ( .gnd!(gnd!), .vdd!(vdd!), .IN0(_2701_), .IN1(PCU_ePC_3_), .Q(_2642__3_), .S(_2643__bF_buf4) );
INX1 INX1_205 ( .gnd!(gnd!), .vdd!(vdd!), .A(PCU_ePC_4_), .Q(_2702_) );
NA2X1 NA2X1_773 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2654_), .B(_2653_), .Q(_2703_) );
NO2I1X1 NO2I1X1_45 ( .gnd!(gnd!), .vdd!(vdd!), .AN(PC1_1_), .B(_2650__bF_buf2), .Q(_2704_) );
AN211X1 AN211X1_15 ( .gnd!(gnd!), .vdd!(vdd!), .A(PC_1_), .B(_2650__bF_buf2), .C(_2663_), .D(_2704_), .Q(_2705_) );
ON21X1 ON21X1_320 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2705_), .B(_2703_), .C(_2665_), .Q(_2706_) );
NA3X1 NA3X1_19 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2672_), .B(_2678_), .C(_2677_), .Q(_2707_) );
ON21X1 ON21X1_321 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2674_), .B(_2673_), .C(_2676_), .Q(_2708_) );
AN22X1 AN22X1_72 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2691_), .B(_2694_), .C(_2707_), .D(_2708_), .Q(_2709_) );
AN21X1 AN21X1_159 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2693_), .B(_2692_), .C(_2688_), .Q(_2710_) );
NA3X1 NA3X1_20 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2688_), .B(_2692_), .C(_2693_), .Q(_2711_) );
NA2X1 NA2X1_774 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2696_), .B(_2711_), .Q(_2712_) );
NA2I1X1 NA2I1X1_114 ( .gnd!(gnd!), .vdd!(vdd!), .AN(_2710_), .B(_2712_), .Q(_2713_) );
AN21X1 AN21X1_160 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2706_), .B(_2709_), .C(_2713_), .Q(_2714_) );
NA2X1 NA2X1_775 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_cu_pc_s2_bF_buf3), .B(I1_4_), .Q(_2715_) );
ON21X1 ON21X1_322 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_cu_pc_s2_bF_buf6), .B(CTRL_cu_pc_s3_bF_buf3), .C(PC1_4_), .Q(_2716_) );
NA2X1 NA2X1_776 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2650__bF_buf2), .B(PC_4_), .Q(_2717_) );
NA3X1 NA3X1_21 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2715_), .B(_2716_), .C(_2717_), .Q(_2718_) );
NA2X1 NA2X1_777 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2717_), .B(_2716_), .Q(_2719_) );
NA2I1X1 NA2I1X1_115 ( .gnd!(gnd!), .vdd!(vdd!), .AN(_2715_), .B(_2719_), .Q(_2720_) );
NA2X1 NA2X1_778 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2720_), .B(_2718_), .Q(_2721_) );
NA2X1 NA2X1_779 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2714_), .B(_2721_), .Q(_2722_) );
AN22X1 AN22X1_73 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_cu_pc_s2_bF_buf3), .B(I1_3_), .C(_2693_), .D(_2692_), .Q(_2723_) );
AN211X1 AN211X1_16 ( .gnd!(gnd!), .vdd!(vdd!), .A(PC_3_), .B(_2650__bF_buf2), .C(_2688_), .D(_2689_), .Q(_2724_) );
ON211X1 ON211X1_112 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2724_), .B(_2723_), .C(_2675_), .D(_2679_), .Q(_2725_) );
AN21X1 AN21X1_161 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2696_), .B(_2711_), .C(_2710_), .Q(_2726_) );
ON21X1 ON21X1_323 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2725_), .B(_2671_), .C(_2726_), .Q(_2727_) );
AN21X1 AN21X1_162 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2717_), .B(_2716_), .C(_2715_), .Q(_2728_) );
NO2I1X1 NO2I1X1_46 ( .gnd!(gnd!), .vdd!(vdd!), .AN(_2718_), .B(_2728_), .Q(_2729_) );
NA2X1 NA2X1_780 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2727_), .B(_2729_), .Q(_2730_) );
AND2X2 AND2X2_81 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2730_), .B(_2686__bF_buf3), .Q(_2731_) );
AO22X2 AO22X2_39 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_IDEC1_cu_jalr_inst_bF_buf5), .B(ALU_r_4_), .C(_2731_), .D(_2722_), .Q(_2732_) );
MU2IX1 MU2IX1_110 ( .gnd!(gnd!), .vdd!(vdd!), .IN0(_2732_), .IN1(PC_4_), .Q(_2733_), .S(_2647__bF_buf1) );
MU2IX1 MU2IX1_111 ( .gnd!(gnd!), .vdd!(vdd!), .IN0(_2733_), .IN1(_2702_), .Q(_2642__4_), .S(_2643__bF_buf1) );
INX1 INX1_206 ( .gnd!(gnd!), .vdd!(vdd!), .A(PCU_ePC_5_), .Q(_2734_) );
NA2X1 NA2X1_781 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2730_), .B(_2720_), .Q(_2735_) );
NA2X1 NA2X1_782 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_cu_pc_s2_bF_buf5), .B(I1_5_), .Q(_2736_) );
ON21X1 ON21X1_324 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_cu_pc_s2_bF_buf6), .B(CTRL_cu_pc_s3_bF_buf0), .C(PC1_5_), .Q(_2737_) );
NA2X1 NA2X1_783 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2650__bF_buf2), .B(PC_5_), .Q(_2738_) );
NA3X1 NA3X1_22 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2736_), .B(_2737_), .C(_2738_), .Q(_2739_) );
NA2X1 NA2X1_784 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2738_), .B(_2737_), .Q(_2740_) );
NA2I1X1 NA2I1X1_116 ( .gnd!(gnd!), .vdd!(vdd!), .AN(_2736_), .B(_2740_), .Q(_2741_) );
NA2X1 NA2X1_785 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2741_), .B(_2739_), .Q(_2742_) );
EN2X1 EN2X1_24 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2735_), .B(_2742_), .Q(_2743_) );
MU2X1 MU2X1_228 ( .gnd!(gnd!), .vdd!(vdd!), .IN0(_2743_), .IN1(ALU_r_5_), .Q(_2744_), .S(CTRL_IDEC1_cu_jalr_inst_bF_buf5) );
MU2IX1 MU2IX1_112 ( .gnd!(gnd!), .vdd!(vdd!), .IN0(_2744_), .IN1(PC_5_), .Q(_2745_), .S(_2647__bF_buf2) );
MU2IX1 MU2IX1_113 ( .gnd!(gnd!), .vdd!(vdd!), .IN0(_2745_), .IN1(_2734_), .Q(_2642__5_), .S(_2643__bF_buf5) );
INX1 INX1_207 ( .gnd!(gnd!), .vdd!(vdd!), .A(PCU_ePC_6_), .Q(_2746_) );
NA2X1 NA2X1_786 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2728_), .B(_2739_), .Q(_2747_) );
NA2X1 NA2X1_787 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2747_), .B(_2741_), .Q(_2748_) );
NO2X1 NO2X1_342 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2721_), .B(_2742_), .Q(_2749_) );
AN21X1 AN21X1_163 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2727_), .B(_2749_), .C(_2748_), .Q(_2750_) );
NA2X1 NA2X1_788 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_cu_pc_s2_bF_buf5), .B(I1_6_), .Q(_2751_) );
OA21X4 OA21X4_3 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_cu_pc_s2_bF_buf5), .B(CTRL_cu_pc_s3_bF_buf0), .C(PC1_6_), .Q(_2752_) );
NO3I1X1 NO3I1X1_5 ( .gnd!(gnd!), .vdd!(vdd!), .AN(PC_6_), .B(CTRL_cu_pc_s2_bF_buf5), .C(CTRL_cu_pc_s3_bF_buf0), .Q(_2753_) );
ON21X1 ON21X1_325 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2752_), .B(_2753_), .C(_2751_), .Q(_2754_) );
ON21X1 ON21X1_326 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_cu_pc_s2_bF_buf5), .B(CTRL_cu_pc_s3_bF_buf0), .C(PC1_6_), .Q(_2755_) );
NA2X1 NA2X1_789 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2650__bF_buf4), .B(PC_6_), .Q(_2756_) );
NA3I1X1 NA3I1X1_118 ( .gnd!(gnd!), .vdd!(vdd!), .AN(_2751_), .B(_2755_), .C(_2756_), .Q(_2757_) );
NA2X1 NA2X1_790 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2754_), .B(_2757_), .Q(_2758_) );
EN2X1 EN2X1_25 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2750_), .B(_2758_), .Q(_2759_) );
MU2X1 MU2X1_229 ( .gnd!(gnd!), .vdd!(vdd!), .IN0(_2759_), .IN1(ALU_r_6_), .Q(_2760_), .S(CTRL_IDEC1_cu_jalr_inst_bF_buf5) );
MU2IX1 MU2IX1_114 ( .gnd!(gnd!), .vdd!(vdd!), .IN0(_2760_), .IN1(PC_6_), .Q(_2761_), .S(_2647__bF_buf2) );
MU2IX1 MU2IX1_115 ( .gnd!(gnd!), .vdd!(vdd!), .IN0(_2761_), .IN1(_2746_), .Q(_2642__6_), .S(_2643__bF_buf5) );
NA2X1 NA2X1_791 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2643__bF_buf0), .B(PCU_ePC_7_), .Q(_2762_) );
AN21X1 AN21X1_164 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2756_), .B(_2755_), .C(_2751_), .Q(_2763_) );
NA2I1X1 NA2I1X1_117 ( .gnd!(gnd!), .vdd!(vdd!), .AN(_2750_), .B(_2758_), .Q(_2764_) );
NA2I1X1 NA2I1X1_118 ( .gnd!(gnd!), .vdd!(vdd!), .AN(_2763_), .B(_2764_), .Q(_2765_) );
AND2X2 AND2X2_82 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_cu_pc_s2_bF_buf5), .B(I1_7_), .Q(_2766_) );
NO2I1X1 NO2I1X1_47 ( .gnd!(gnd!), .vdd!(vdd!), .AN(PC1_7_), .B(_2650__bF_buf4), .Q(_2767_) );
NO3I1X1 NO3I1X1_6 ( .gnd!(gnd!), .vdd!(vdd!), .AN(PC_7_), .B(CTRL_cu_pc_s2_bF_buf4), .C(CTRL_cu_pc_s3_bF_buf2), .Q(_2768_) );
ON21X1 ON21X1_327 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2767_), .B(_2768_), .C(_2766_), .Q(_2769_) );
NA2X1 NA2X1_792 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_cu_pc_s2_bF_buf5), .B(I1_7_), .Q(_2770_) );
ON21X1 ON21X1_328 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_cu_pc_s2_bF_buf5), .B(CTRL_cu_pc_s3_bF_buf0), .C(PC1_7_), .Q(_2771_) );
NA2X1 NA2X1_793 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2650__bF_buf4), .B(PC_7_), .Q(_2772_) );
NA3X1 NA3X1_23 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2770_), .B(_2771_), .C(_2772_), .Q(_2773_) );
NA2X1 NA2X1_794 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2769_), .B(_2773_), .Q(_2774_) );
EN2X1 EN2X1_26 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2765_), .B(_2774_), .Q(_2775_) );
MU2X1 MU2X1_230 ( .gnd!(gnd!), .vdd!(vdd!), .IN0(_2775_), .IN1(ALU_r_7_), .Q(_2776_), .S(CTRL_IDEC1_cu_jalr_inst_bF_buf5) );
NO2X1 NO2X1_343 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2647__bF_buf0), .B(_2776_), .Q(_2777_) );
NO2X1 NO2X1_344 ( .gnd!(gnd!), .vdd!(vdd!), .A(PC_7_), .B(_2646__bF_buf1), .Q(_2778_) );
ON31X1 ON31X1_87 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2643__bF_buf0), .B(_2778_), .C(_2777_), .D(_2762_), .Q(_2642__7_) );
AN21X1 AN21X1_165 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2738_), .B(_2737_), .C(_2736_), .Q(_2779_) );
NO2I1X1 NO2I1X1_48 ( .gnd!(gnd!), .vdd!(vdd!), .AN(_2739_), .B(_2779_), .Q(_2780_) );
ON21X1 ON21X1_329 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2767_), .B(_2768_), .C(_2770_), .Q(_2781_) );
NA3I1X1 NA3I1X1_119 ( .gnd!(gnd!), .vdd!(vdd!), .AN(_2770_), .B(_2771_), .C(_2772_), .Q(_2782_) );
AN22X1 AN22X1_74 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2754_), .B(_2757_), .C(_2781_), .D(_2782_), .Q(_2783_) );
NA3X1 NA3X1_24 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2783_), .B(_2729_), .C(_2780_), .Q(_2784_) );
NA2X1 NA2X1_795 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2763_), .B(_2773_), .Q(_2785_) );
NA2X1 NA2X1_796 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2785_), .B(_2769_), .Q(_2786_) );
AN21X1 AN21X1_166 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2748_), .B(_2783_), .C(_2786_), .Q(_2787_) );
ON21X1 ON21X1_330 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2714_), .B(_2784_), .C(_2787_), .Q(_2788_) );
NA2X1 NA2X1_797 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_cu_pc_s2_bF_buf6), .B(I1_8_), .Q(_2789_) );
ON21X1 ON21X1_331 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_cu_pc_s2_bF_buf2), .B(CTRL_cu_pc_s3_bF_buf4), .C(PC1_8_), .Q(_2790_) );
NA2X1 NA2X1_798 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2650__bF_buf1), .B(PC_8_), .Q(_2791_) );
NA2X1 NA2X1_799 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2791_), .B(_2790_), .Q(_2792_) );
NA2X1 NA2X1_800 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2792_), .B(_2789_), .Q(_2793_) );
NA3I1X1 NA3I1X1_120 ( .gnd!(gnd!), .vdd!(vdd!), .AN(_2789_), .B(_2790_), .C(_2791_), .Q(_2794_) );
NA2X1 NA2X1_801 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2793_), .B(_2794_), .Q(_2795_) );
NO2X1 NO2X1_345 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2795_), .B(_2788_), .Q(_2796_) );
AND2X2 AND2X2_83 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2788_), .B(_2795_), .Q(_2797_) );
NA2X1 NA2X1_802 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_IDEC1_cu_jalr_inst_bF_buf4), .B(ALU_r_8_), .Q(_2798_) );
ON31X1 ON31X1_88 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_IDEC1_cu_jalr_inst_bF_buf1), .B(_2796_), .C(_2797_), .D(_2798_), .Q(_2799_) );
MU2X1 MU2X1_231 ( .gnd!(gnd!), .vdd!(vdd!), .IN0(_2799_), .IN1(PC_8_), .Q(_2800_), .S(_2647__bF_buf4) );
MU2X1 MU2X1_232 ( .gnd!(gnd!), .vdd!(vdd!), .IN0(_2800_), .IN1(PCU_ePC_8_), .Q(_2642__8_), .S(_2643__bF_buf4) );
NA2X1 NA2X1_803 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_IDEC1_cu_jalr_inst_bF_buf4), .B(ALU_r_9_), .Q(_2801_) );
NA2I1X1 NA2I1X1_119 ( .gnd!(gnd!), .vdd!(vdd!), .AN(_2789_), .B(_2792_), .Q(_2802_) );
NA2X1 NA2X1_804 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_cu_pc_s2_bF_buf3), .B(I1_9_), .Q(_2803_) );
ON21X1 ON21X1_332 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_cu_pc_s2_bF_buf6), .B(CTRL_cu_pc_s3_bF_buf1), .C(PC1_9_), .Q(_2804_) );
NA2X1 NA2X1_805 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2650__bF_buf1), .B(PC_9_), .Q(_2805_) );
AN21X1 AN21X1_167 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2805_), .B(_2804_), .C(_2803_), .Q(_2806_) );
INX1 INX1_208 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2803_), .Q(_2807_) );
NA2X1 NA2X1_806 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2805_), .B(_2804_), .Q(_2808_) );
NO2X1 NO2X1_346 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2807_), .B(_2808_), .Q(_2809_) );
AN211X1 AN211X1_17 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2794_), .B(_2793_), .C(_2806_), .D(_2809_), .Q(_2810_) );
NA2X1 NA2X1_807 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2788_), .B(_2810_), .Q(_2811_) );
ON31X1 ON31X1_89 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2802_), .B(_2806_), .C(_2809_), .D(_2811_), .Q(_2812_) );
AN21X1 AN21X1_168 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2791_), .B(_2790_), .C(_2789_), .Q(_2813_) );
NA2X1 NA2X1_808 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2808_), .B(_2807_), .Q(_2814_) );
NA3X1 NA3X1_25 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2803_), .B(_2804_), .C(_2805_), .Q(_2815_) );
AN211X1 AN211X1_18 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2814_), .B(_2815_), .C(_2813_), .D(_2797_), .Q(_2816_) );
ON31X1 ON31X1_90 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_IDEC1_cu_jalr_inst_bF_buf0), .B(_2812_), .C(_2816_), .D(_2801_), .Q(_2817_) );
MU2X1 MU2X1_233 ( .gnd!(gnd!), .vdd!(vdd!), .IN0(_2817_), .IN1(PC_9_), .Q(_2818_), .S(_2647__bF_buf2) );
MU2X1 MU2X1_234 ( .gnd!(gnd!), .vdd!(vdd!), .IN0(_2818_), .IN1(PCU_ePC_9_), .Q(_2642__9_), .S(_2643__bF_buf5) );
NA2X1 NA2X1_809 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2643__bF_buf4), .B(PCU_ePC_10_), .Q(_2819_) );
AN21X1 AN21X1_169 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2813_), .B(_2815_), .C(_2806_), .Q(_2820_) );
NA2X1 NA2X1_810 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2811_), .B(_2820_), .Q(_2821_) );
NA2X1 NA2X1_811 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_cu_pc_s2_bF_buf7), .B(I1_10_), .Q(_2822_) );
NO2I1X1 NO2I1X1_49 ( .gnd!(gnd!), .vdd!(vdd!), .AN(PC1_10_), .B(_2650__bF_buf4), .Q(_2823_) );
NO3I1X1 NO3I1X1_7 ( .gnd!(gnd!), .vdd!(vdd!), .AN(PC_10_), .B(CTRL_cu_pc_s2_bF_buf7), .C(CTRL_cu_pc_s3_bF_buf4), .Q(_2824_) );
ON21X1 ON21X1_333 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2823_), .B(_2824_), .C(_2822_), .Q(_2825_) );
ON21X1 ON21X1_334 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_cu_pc_s2_bF_buf7), .B(CTRL_cu_pc_s3_bF_buf4), .C(PC1_10_), .Q(_2826_) );
NA2X1 NA2X1_812 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2650__bF_buf1), .B(PC_10_), .Q(_2827_) );
NA3I1X1 NA3I1X1_121 ( .gnd!(gnd!), .vdd!(vdd!), .AN(_2822_), .B(_2826_), .C(_2827_), .Q(_2828_) );
NA2X1 NA2X1_813 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2825_), .B(_2828_), .Q(_2829_) );
NA2X1 NA2X1_814 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2821_), .B(_2829_), .Q(_2830_) );
OR2X2 OR2X2_24 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2821_), .B(_2829_), .Q(_2831_) );
NA2X1 NA2X1_815 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2831_), .B(_2830_), .Q(_2832_) );
NA2X1 NA2X1_816 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2832_), .B(_2686__bF_buf2), .Q(_2833_) );
NA2I1X1 NA2I1X1_120 ( .gnd!(gnd!), .vdd!(vdd!), .AN(ALU_r_10_), .B(CTRL_IDEC1_cu_jalr_inst_bF_buf1), .Q(_2834_) );
INX1 INX1_209 ( .gnd!(gnd!), .vdd!(vdd!), .A(PC_10_), .Q(_2835_) );
NO2X1 NO2X1_347 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2835_), .B(_2646__bF_buf3), .Q(_2836_) );
AN31X1 AN31X1_79 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2646__bF_buf3), .B(_2834_), .C(_2833_), .D(_2836_), .Q(_2837_) );
ON21X1 ON21X1_335 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2837_), .B(_2643__bF_buf4), .C(_2819_), .Q(_2642__10_) );
NO2X1 NO2X1_348 ( .gnd!(gnd!), .vdd!(vdd!), .A(ALU_r_11_), .B(_2686__bF_buf2), .Q(_2838_) );
AN21X1 AN21X1_170 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2827_), .B(_2826_), .C(_2822_), .Q(_2839_) );
NA2X1 NA2X1_817 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_cu_pc_s2_bF_buf3), .B(I1_11_), .Q(_2840_) );
NO2I1X1 NO2I1X1_50 ( .gnd!(gnd!), .vdd!(vdd!), .AN(PC1_11_), .B(_2650__bF_buf1), .Q(_2841_) );
NO3I1X1 NO3I1X1_8 ( .gnd!(gnd!), .vdd!(vdd!), .AN(PC_11_), .B(CTRL_cu_pc_s2_bF_buf7), .C(CTRL_cu_pc_s3_bF_buf4), .Q(_2842_) );
ON21X1 ON21X1_336 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2841_), .B(_2842_), .C(_2840_), .Q(_2843_) );
NA2I1X1 NA2I1X1_121 ( .gnd!(gnd!), .vdd!(vdd!), .AN(_2650__bF_buf1), .B(PC1_11_), .Q(_2844_) );
NA2X1 NA2X1_818 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2650__bF_buf1), .B(PC_11_), .Q(_2845_) );
NA3I1X1 NA3I1X1_122 ( .gnd!(gnd!), .vdd!(vdd!), .AN(_2840_), .B(_2845_), .C(_2844_), .Q(_2846_) );
NA2X1 NA2X1_819 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2846_), .B(_2843_), .Q(_2847_) );
NA3I1X1 NA3I1X1_123 ( .gnd!(gnd!), .vdd!(vdd!), .AN(_2839_), .B(_2847_), .C(_2830_), .Q(_2848_) );
ON211X1 ON211X1_113 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2823_), .B(_2824_), .C(CTRL_cu_pc_s2_bF_buf7), .D(I1_10_), .Q(_2849_) );
AND2X2 AND2X2_84 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_cu_pc_s2_bF_buf3), .B(I1_11_), .Q(_2850_) );
ON21X1 ON21X1_337 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2841_), .B(_2842_), .C(_2850_), .Q(_2851_) );
INX1 INX1_210 ( .gnd!(gnd!), .vdd!(vdd!), .A(PC1_11_), .Q(_2852_) );
ON211X1 ON211X1_114 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2852_), .B(_2650__bF_buf1), .C(_2845_), .D(_2840_), .Q(_2853_) );
AO22X2 AO22X2_40 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2851_), .B(_2853_), .C(_2830_), .D(_2849_), .Q(_2854_) );
AN31X1 AN31X1_80 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2686__bF_buf2), .B(_2848_), .C(_2854_), .D(_2838_), .Q(_2855_) );
MU2X1 MU2X1_235 ( .gnd!(gnd!), .vdd!(vdd!), .IN0(_2855_), .IN1(PC_11_), .Q(_2856_), .S(_2647__bF_buf0) );
MU2X1 MU2X1_236 ( .gnd!(gnd!), .vdd!(vdd!), .IN0(_2856_), .IN1(PCU_ePC_11_), .Q(_2642__11_), .S(_2643__bF_buf5) );
NA2X1 NA2X1_820 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_IDEC1_cu_jalr_inst_bF_buf1), .B(ALU_r_12_), .Q(_2857_) );
AN21X1 AN21X1_171 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2728_), .B(_2739_), .C(_2779_), .Q(_2858_) );
AN22X1 AN22X1_75 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_cu_pc_s2_bF_buf5), .B(I1_6_), .C(_2756_), .D(_2755_), .Q(_2859_) );
AN211X1 AN211X1_19 ( .gnd!(gnd!), .vdd!(vdd!), .A(PC_6_), .B(_2650__bF_buf4), .C(_2751_), .D(_2752_), .Q(_2860_) );
ON211X1 ON211X1_115 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2860_), .B(_2859_), .C(_2769_), .D(_2773_), .Q(_2861_) );
AN21X1 AN21X1_172 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2772_), .B(_2771_), .C(_2770_), .Q(_2862_) );
AN21X1 AN21X1_173 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2763_), .B(_2773_), .C(_2862_), .Q(_2863_) );
ON21X1 ON21X1_338 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2861_), .B(_2858_), .C(_2863_), .Q(_2864_) );
AN31X1 AN31X1_81 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2749_), .B(_2783_), .C(_2727_), .D(_2864_), .Q(_2865_) );
AN22X1 AN22X1_76 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2825_), .B(_2828_), .C(_2843_), .D(_2846_), .Q(_2866_) );
NA2X1 NA2X1_821 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2810_), .B(_2866_), .Q(_2867_) );
ON21X1 ON21X1_339 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2809_), .B(_2802_), .C(_2814_), .Q(_2868_) );
NA2X1 NA2X1_822 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2849_), .B(_2851_), .Q(_2869_) );
AN22X1 AN22X1_77 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2853_), .B(_2869_), .C(_2868_), .D(_2866_), .Q(_2870_) );
ON21X1 ON21X1_340 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2865_), .B(_2867_), .C(_2870_), .Q(_2871_) );
NA2X1 NA2X1_823 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_cu_pc_s2_bF_buf0), .B(I1_12_), .Q(_2872_) );
NO2I1X1 NO2I1X1_51 ( .gnd!(gnd!), .vdd!(vdd!), .AN(PC1_12_), .B(_2650__bF_buf4), .Q(_2873_) );
NO3I1X1 NO3I1X1_9 ( .gnd!(gnd!), .vdd!(vdd!), .AN(PC_12_), .B(CTRL_cu_pc_s2_bF_buf0), .C(CTRL_cu_pc_s3_bF_buf2), .Q(_2874_) );
ON21X1 ON21X1_341 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2873_), .B(_2874_), .C(_2872_), .Q(_2875_) );
INX1 INX1_211 ( .gnd!(gnd!), .vdd!(vdd!), .A(PC1_12_), .Q(_2876_) );
AND2X2 AND2X2_85 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_cu_pc_s2_bF_buf0), .B(I1_12_), .Q(_2877_) );
NA2X1 NA2X1_824 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2650__bF_buf3), .B(PC_12_), .Q(_2878_) );
ON211X1 ON211X1_116 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2876_), .B(_2650__bF_buf3), .C(_2878_), .D(_2877_), .Q(_2879_) );
NA2X1 NA2X1_825 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2879_), .B(_2875_), .Q(_2880_) );
NA2X1 NA2X1_826 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2871_), .B(_2880_), .Q(_2881_) );
NO2X1 NO2X1_349 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2880_), .B(_2871_), .Q(_2882_) );
NA3I1X1 NA3I1X1_124 ( .gnd!(gnd!), .vdd!(vdd!), .AN(_2882_), .B(_2686__bF_buf0), .C(_2881_), .Q(_2883_) );
NA2X1 NA2X1_827 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2883_), .B(_2857_), .Q(_2884_) );
MU2X1 MU2X1_237 ( .gnd!(gnd!), .vdd!(vdd!), .IN0(_2884_), .IN1(PC_12_), .Q(_2885_), .S(_2647__bF_buf1) );
MU2X1 MU2X1_238 ( .gnd!(gnd!), .vdd!(vdd!), .IN0(_2885_), .IN1(PCU_ePC_12_), .Q(_2642__12_), .S(_2643__bF_buf1) );
NA2X1 NA2X1_828 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_IDEC1_cu_jalr_inst_bF_buf2), .B(ALU_r_13_), .Q(_2886_) );
ON21X1 ON21X1_342 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2873_), .B(_2874_), .C(_2877_), .Q(_2887_) );
NA2X1 NA2X1_829 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_cu_pc_s2_bF_buf0), .B(I1_13_), .Q(_2888_) );
INX1 INX1_212 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2888_), .Q(_2889_) );
ON21X1 ON21X1_343 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_cu_pc_s2_bF_buf0), .B(CTRL_cu_pc_s3_bF_buf2), .C(PC1_13_), .Q(_2890_) );
NA2X1 NA2X1_830 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2650__bF_buf3), .B(PC_13_), .Q(_2891_) );
NA2X1 NA2X1_831 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2891_), .B(_2890_), .Q(_2892_) );
NA2X1 NA2X1_832 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2892_), .B(_2889_), .Q(_2893_) );
NA3X1 NA3X1_26 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2888_), .B(_2890_), .C(_2891_), .Q(_2894_) );
NA2X1 NA2X1_833 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2893_), .B(_2894_), .Q(_2895_) );
AND3X4 AND3X4_15 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2881_), .B(_2887_), .C(_2895_), .Q(_2896_) );
AN21X1 AN21X1_174 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2891_), .B(_2890_), .C(_2888_), .Q(_2897_) );
NO2X1 NO2X1_350 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2889_), .B(_2892_), .Q(_2898_) );
ON31X1 ON31X1_91 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2887_), .B(_2897_), .C(_2898_), .D(_2686__bF_buf0), .Q(_2899_) );
NO2X1 NO2X1_351 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2895_), .B(_2881_), .Q(_2900_) );
ON31X1 ON31X1_92 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2899_), .B(_2900_), .C(_2896_), .D(_2886_), .Q(_2901_) );
MU2X1 MU2X1_239 ( .gnd!(gnd!), .vdd!(vdd!), .IN0(_2901_), .IN1(PC_13_), .Q(_2902_), .S(_2647__bF_buf0) );
MU2X1 MU2X1_240 ( .gnd!(gnd!), .vdd!(vdd!), .IN0(_2902_), .IN1(PCU_ePC_13_), .Q(_2642__13_), .S(_2643__bF_buf1) );
NA2X1 NA2X1_834 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2643__bF_buf2), .B(PCU_ePC_14_), .Q(_2903_) );
AND2X2 AND2X2_86 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_IDEC1_cu_jalr_inst_bF_buf4), .B(ALU_r_14_), .Q(_2904_) );
ON21X1 ON21X1_344 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2898_), .B(_2887_), .C(_2893_), .Q(_2905_) );
NO2X1 NO2X1_352 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2905_), .B(_2900_), .Q(_2906_) );
NO2I1X1 NO2I1X1_52 ( .gnd!(gnd!), .vdd!(vdd!), .AN(PC1_14_), .B(_2650__bF_buf4), .Q(_2907_) );
NO3I1X1 NO3I1X1_10 ( .gnd!(gnd!), .vdd!(vdd!), .AN(PC_14_), .B(CTRL_cu_pc_s2_bF_buf4), .C(CTRL_cu_pc_s3_bF_buf4), .Q(_2908_) );
AN211X1 AN211X1_20 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_cu_pc_s2_bF_buf4), .B(I1_14_), .C(_2908_), .D(_2907_), .Q(_2909_) );
INX1 INX1_213 ( .gnd!(gnd!), .vdd!(vdd!), .A(PC_14_), .Q(_2910_) );
NA2X1 NA2X1_835 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_cu_pc_s2_bF_buf4), .B(I1_14_), .Q(_2911_) );
NO2X1 NO2X1_353 ( .gnd!(gnd!), .vdd!(vdd!), .A(PC1_14_), .B(_2650__bF_buf7), .Q(_2912_) );
AN211X1 AN211X1_21 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2910_), .B(_2650__bF_buf7), .C(_2911_), .D(_2912_), .Q(_2913_) );
NO2X1 NO2X1_354 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2913_), .B(_2909_), .Q(_2914_) );
INX1 INX1_214 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2914_), .Q(_2915_) );
NA2X1 NA2X1_836 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2906_), .B(_2915_), .Q(_2916_) );
NA2I1X1 NA2I1X1_122 ( .gnd!(gnd!), .vdd!(vdd!), .AN(_2906_), .B(_2914_), .Q(_2917_) );
AND3X4 AND3X4_16 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2917_), .B(_2686__bF_buf0), .C(_2916_), .Q(_2918_) );
NO3X1 NO3X1_19 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2918_), .B(_2647__bF_buf3), .C(_2904_), .Q(_2919_) );
ON21X1 ON21X1_345 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2646__bF_buf2), .B(PC_14_), .C(CTRL_cu_ld_epc), .Q(_2920_) );
ON21X1 ON21X1_346 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2919_), .B(_2920_), .C(_2903_), .Q(_2642__14_) );
NA2X1 NA2X1_837 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2643__bF_buf1), .B(PCU_ePC_15_), .Q(_2921_) );
NO2X1 NO2X1_355 ( .gnd!(gnd!), .vdd!(vdd!), .A(ALU_r_15_), .B(_2686__bF_buf0), .Q(_2922_) );
ON211X1 ON211X1_117 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2907_), .B(_2908_), .C(CTRL_cu_pc_s2_bF_buf4), .D(I1_14_), .Q(_2923_) );
ON21X1 ON21X1_347 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2906_), .B(_2915_), .C(_2923_), .Q(_2924_) );
NA2X1 NA2X1_838 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_cu_pc_s2_bF_buf0), .B(I1_15_), .Q(_2925_) );
ON21X1 ON21X1_348 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_cu_pc_s2_bF_buf0), .B(CTRL_cu_pc_s3_bF_buf2), .C(PC1_15_), .Q(_2926_) );
NA2X1 NA2X1_839 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2650__bF_buf3), .B(PC_15_), .Q(_2927_) );
AN21X1 AN21X1_175 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2927_), .B(_2926_), .C(_2925_), .Q(_2928_) );
NA3X1 NA3X1_27 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2925_), .B(_2926_), .C(_2927_), .Q(_2929_) );
NO2I1X1 NO2I1X1_53 ( .gnd!(gnd!), .vdd!(vdd!), .AN(_2929_), .B(_2928_), .Q(_2930_) );
NA2I1X1 NA2I1X1_123 ( .gnd!(gnd!), .vdd!(vdd!), .AN(_2930_), .B(_2924_), .Q(_2931_) );
NA3I1X1 NA3I1X1_125 ( .gnd!(gnd!), .vdd!(vdd!), .AN(_2913_), .B(_2930_), .C(_2917_), .Q(_2932_) );
AN31X1 AN31X1_82 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2686__bF_buf0), .B(_2931_), .C(_2932_), .D(_2922_), .Q(_2933_) );
INX1 INX1_215 ( .gnd!(gnd!), .vdd!(vdd!), .A(PC_15_), .Q(_2934_) );
NA2X1 NA2X1_840 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2647__bF_buf1), .B(_2934_), .Q(_2935_) );
ON211X1 ON211X1_118 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2933_), .B(_2647__bF_buf2), .C(CTRL_cu_ld_epc), .D(_2935_), .Q(_2936_) );
NA2X1 NA2X1_841 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2936_), .B(_2921_), .Q(_2642__15_) );
AN22X1 AN22X1_78 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_cu_pc_s2_bF_buf7), .B(I1_10_), .C(_2827_), .D(_2826_), .Q(_2937_) );
NO3X1 NO3X1_20 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2823_), .B(_2824_), .C(_2822_), .Q(_2938_) );
ON211X1 ON211X1_119 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2938_), .B(_2937_), .C(_2851_), .D(_2853_), .Q(_2939_) );
ON211X1 ON211X1_120 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2876_), .B(_2650__bF_buf3), .C(_2878_), .D(_2872_), .Q(_2940_) );
AN22X1 AN22X1_79 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_cu_pc_s2_bF_buf0), .B(I1_13_), .C(_2891_), .D(_2890_), .Q(_2941_) );
NO2I1X1 NO2I1X1_54 ( .gnd!(gnd!), .vdd!(vdd!), .AN(PC1_13_), .B(_2650__bF_buf4), .Q(_2942_) );
AN211X1 AN211X1_22 ( .gnd!(gnd!), .vdd!(vdd!), .A(PC_13_), .B(_2650__bF_buf3), .C(_2888_), .D(_2942_), .Q(_2943_) );
ON211X1 ON211X1_121 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2943_), .B(_2941_), .C(_2887_), .D(_2940_), .Q(_2944_) );
INX1 INX1_216 ( .gnd!(gnd!), .vdd!(vdd!), .A(PC1_14_), .Q(_2945_) );
NA2X1 NA2X1_842 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2650__bF_buf7), .B(PC_14_), .Q(_2946_) );
ON211X1 ON211X1_122 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2945_), .B(_2650__bF_buf3), .C(_2946_), .D(_2911_), .Q(_2947_) );
AN22X1 AN22X1_80 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_cu_pc_s2_bF_buf0), .B(I1_15_), .C(_2927_), .D(_2926_), .Q(_2948_) );
NO2I1X1 NO2I1X1_55 ( .gnd!(gnd!), .vdd!(vdd!), .AN(PC1_15_), .B(_2650__bF_buf4), .Q(_2949_) );
AN211X1 AN211X1_23 ( .gnd!(gnd!), .vdd!(vdd!), .A(PC_15_), .B(_2650__bF_buf3), .C(_2925_), .D(_2949_), .Q(_2950_) );
ON211X1 ON211X1_123 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2950_), .B(_2948_), .C(_2947_), .D(_2923_), .Q(_2951_) );
NO2X1 NO2X1_356 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2944_), .B(_2951_), .Q(_2952_) );
NA3I1X1 NA3I1X1_126 ( .gnd!(gnd!), .vdd!(vdd!), .AN(_2939_), .B(_2810_), .C(_2952_), .Q(_2953_) );
NA2X1 NA2X1_843 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2869_), .B(_2853_), .Q(_2954_) );
ON21X1 ON21X1_349 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2939_), .B(_2820_), .C(_2954_), .Q(_2955_) );
NA2I1X1 NA2I1X1_124 ( .gnd!(gnd!), .vdd!(vdd!), .AN(_2873_), .B(_2878_), .Q(_2956_) );
AN31X1 AN31X1_83 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2877_), .B(_2894_), .C(_2956_), .D(_2897_), .Q(_2957_) );
AN21X1 AN21X1_176 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2913_), .B(_2929_), .C(_2928_), .Q(_2958_) );
ON21X1 ON21X1_350 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2957_), .B(_2951_), .C(_2958_), .Q(_2959_) );
AN21X1 AN21X1_177 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2952_), .B(_2955_), .C(_2959_), .Q(_2960_) );
ON21X1 ON21X1_351 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2865_), .B(_2953_), .C(_2960_), .Q(_2961_) );
INX1 INX1_217 ( .gnd!(gnd!), .vdd!(vdd!), .A(PC_16_), .Q(_2962_) );
NA2X1 NA2X1_844 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_cu_pc_s2_bF_buf3), .B(I1_16_), .Q(_2963_) );
NO2X1 NO2X1_357 ( .gnd!(gnd!), .vdd!(vdd!), .A(PC1_16_), .B(_2650__bF_buf5), .Q(_2964_) );
AO211X4 AO211X4_1 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2962_), .B(_2650__bF_buf5), .C(_2963_), .D(_2964_), .Q(_2965_) );
MU2IX1 MU2IX1_116 ( .gnd!(gnd!), .vdd!(vdd!), .IN0(PC1_16_), .IN1(PC_16_), .Q(_2966_), .S(_2650__bF_buf5) );
NA2X1 NA2X1_845 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2966_), .B(_2963_), .Q(_2967_) );
NA2X1 NA2X1_846 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2967_), .B(_2965_), .Q(_2968_) );
INX1 INX1_218 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2968_), .Q(_2969_) );
NA2X1 NA2X1_847 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2961_), .B(_2969_), .Q(_2970_) );
NA2X1 NA2X1_848 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2892_), .B(_2888_), .Q(_2971_) );
NA3I1X1 NA3I1X1_127 ( .gnd!(gnd!), .vdd!(vdd!), .AN(_2888_), .B(_2890_), .C(_2891_), .Q(_2972_) );
AN22X1 AN22X1_81 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2879_), .B(_2875_), .C(_2971_), .D(_2972_), .Q(_2973_) );
NA3X1 NA3X1_28 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2930_), .B(_2914_), .C(_2973_), .Q(_2974_) );
NO2X1 NO2X1_358 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2974_), .B(_2867_), .Q(_2975_) );
ON21X1 ON21X1_352 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2945_), .B(_2650__bF_buf7), .C(_2946_), .Q(_2976_) );
NA3I1X1 NA3I1X1_128 ( .gnd!(gnd!), .vdd!(vdd!), .AN(_2911_), .B(_2929_), .C(_2976_), .Q(_2977_) );
NA2I1X1 NA2I1X1_125 ( .gnd!(gnd!), .vdd!(vdd!), .AN(_2928_), .B(_2977_), .Q(_2978_) );
AN31X1 AN31X1_84 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2930_), .B(_2914_), .C(_2905_), .D(_2978_), .Q(_2979_) );
ON21X1 ON21X1_353 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2870_), .B(_2974_), .C(_2979_), .Q(_2980_) );
AN21X1 AN21X1_178 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2788_), .B(_2975_), .C(_2980_), .Q(_2981_) );
NA2X1 NA2X1_849 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2981_), .B(_2968_), .Q(_2982_) );
AND2X2 AND2X2_87 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_IDEC1_cu_jalr_inst_bF_buf2), .B(ALU_r_16_), .Q(_2983_) );
AO31X1 AO31X1_1 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2686__bF_buf1), .B(_2970_), .C(_2982_), .D(_2983_), .Q(_2984_) );
MU2X1 MU2X1_241 ( .gnd!(gnd!), .vdd!(vdd!), .IN0(_2984_), .IN1(PC_16_), .Q(_2985_), .S(_2647__bF_buf4) );
MU2X1 MU2X1_242 ( .gnd!(gnd!), .vdd!(vdd!), .IN0(_2985_), .IN1(PCU_ePC_16_), .Q(_2642__16_), .S(_2643__bF_buf3) );
NA2X1 NA2X1_850 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_cu_pc_s2_bF_buf4), .B(I1_17_), .Q(_2986_) );
INX1 INX1_219 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2986_), .Q(_2987_) );
MU2X1 MU2X1_243 ( .gnd!(gnd!), .vdd!(vdd!), .IN0(PC1_17_), .IN1(PC_17_), .Q(_2988_), .S(_2650__bF_buf7) );
NA2X1 NA2X1_851 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2988_), .B(_2987_), .Q(_2989_) );
MU2IX1 MU2IX1_117 ( .gnd!(gnd!), .vdd!(vdd!), .IN0(PC1_17_), .IN1(PC_17_), .Q(_2990_), .S(_2650__bF_buf7) );
NA2X1 NA2X1_852 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2990_), .B(_2986_), .Q(_2991_) );
NA2X1 NA2X1_853 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2989_), .B(_2991_), .Q(_2992_) );
INX1 INX1_220 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2992_), .Q(_2993_) );
NA2X1 NA2X1_854 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2970_), .B(_2965_), .Q(_2994_) );
NA2X1 NA2X1_855 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2994_), .B(_2993_), .Q(_2995_) );
AN31X1 AN31X1_85 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2965_), .B(_2992_), .C(_2970_), .D(CTRL_IDEC1_cu_jalr_inst_bF_buf2), .Q(_2996_) );
AO22X2 AO22X2_41 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_IDEC1_cu_jalr_inst_bF_buf2), .B(ALU_r_17_), .C(_2995_), .D(_2996_), .Q(_2997_) );
MU2X1 MU2X1_244 ( .gnd!(gnd!), .vdd!(vdd!), .IN0(_2997_), .IN1(PC_17_), .Q(_2998_), .S(_2647__bF_buf0) );
MU2X1 MU2X1_245 ( .gnd!(gnd!), .vdd!(vdd!), .IN0(_2998_), .IN1(PCU_ePC_17_), .Q(_2642__17_), .S(_2643__bF_buf0) );
NA2X1 NA2X1_856 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2643__bF_buf3), .B(PCU_ePC_18_), .Q(_2999_) );
AND2X2 AND2X2_88 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_IDEC1_cu_jalr_inst_bF_buf1), .B(ALU_r_18_), .Q(_3000_) );
NO2X1 NO2X1_359 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2968_), .B(_2992_), .Q(_3001_) );
NO2X1 NO2X1_360 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2987_), .B(_2988_), .Q(_3002_) );
ON21X1 ON21X1_354 ( .gnd!(gnd!), .vdd!(vdd!), .A(_3002_), .B(_2965_), .C(_2989_), .Q(_3003_) );
AN21X1 AN21X1_179 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2961_), .B(_3001_), .C(_3003_), .Q(_3004_) );
NA2X1 NA2X1_857 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_cu_pc_s2_bF_buf3), .B(I1_18_), .Q(_3005_) );
MU2IX1 MU2IX1_118 ( .gnd!(gnd!), .vdd!(vdd!), .IN0(PC1_18_), .IN1(PC_18_), .Q(_3006_), .S(_2650__bF_buf5) );
NA2X1 NA2X1_858 ( .gnd!(gnd!), .vdd!(vdd!), .A(_3006_), .B(_3005_), .Q(_3007_) );
INX1 INX1_221 ( .gnd!(gnd!), .vdd!(vdd!), .A(PC_18_), .Q(_3008_) );
NO2X1 NO2X1_361 ( .gnd!(gnd!), .vdd!(vdd!), .A(PC1_18_), .B(_2650__bF_buf5), .Q(_3009_) );
AO211X4 AO211X4_2 ( .gnd!(gnd!), .vdd!(vdd!), .A(_3008_), .B(_2650__bF_buf0), .C(_3005_), .D(_3009_), .Q(_3010_) );
NA2X1 NA2X1_859 ( .gnd!(gnd!), .vdd!(vdd!), .A(_3007_), .B(_3010_), .Q(_3011_) );
EN2X1 EN2X1_27 ( .gnd!(gnd!), .vdd!(vdd!), .A(_3004_), .B(_3011_), .Q(_3012_) );
NO2X1 NO2X1_362 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_IDEC1_cu_jalr_inst_bF_buf1), .B(_3012_), .Q(_3013_) );
NO3X1 NO3X1_21 ( .gnd!(gnd!), .vdd!(vdd!), .A(_3013_), .B(_2647__bF_buf4), .C(_3000_), .Q(_3014_) );
NO2X1 NO2X1_363 ( .gnd!(gnd!), .vdd!(vdd!), .A(PC_18_), .B(_2646__bF_buf3), .Q(_3015_) );
ON31X1 ON31X1_93 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2643__bF_buf3), .B(_3015_), .C(_3014_), .D(_2999_), .Q(_2642__18_) );
INX1 INX1_222 ( .gnd!(gnd!), .vdd!(vdd!), .A(PC_19_), .Q(_3016_) );
ON21X1 ON21X1_355 ( .gnd!(gnd!), .vdd!(vdd!), .A(_3004_), .B(_3011_), .C(_3010_), .Q(_3017_) );
NA2X1 NA2X1_860 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_cu_pc_s2_bF_buf7), .B(I1_19_), .Q(_3018_) );
INX1 INX1_223 ( .gnd!(gnd!), .vdd!(vdd!), .A(_3018_), .Q(_3019_) );
NO2X1 NO2X1_364 ( .gnd!(gnd!), .vdd!(vdd!), .A(PC1_19_), .B(_2650__bF_buf7), .Q(_3020_) );
AN21X1 AN21X1_180 ( .gnd!(gnd!), .vdd!(vdd!), .A(_3016_), .B(_2650__bF_buf0), .C(_3020_), .Q(_3021_) );
NA2X1 NA2X1_861 ( .gnd!(gnd!), .vdd!(vdd!), .A(_3021_), .B(_3019_), .Q(_3022_) );
MU2IX1 MU2IX1_119 ( .gnd!(gnd!), .vdd!(vdd!), .IN0(PC1_19_), .IN1(PC_19_), .Q(_3023_), .S(_2650__bF_buf7) );
NA2X1 NA2X1_862 ( .gnd!(gnd!), .vdd!(vdd!), .A(_3023_), .B(_3018_), .Q(_3024_) );
AND2X2 AND2X2_89 ( .gnd!(gnd!), .vdd!(vdd!), .A(_3024_), .B(_3022_), .Q(_3025_) );
NA2X1 NA2X1_863 ( .gnd!(gnd!), .vdd!(vdd!), .A(_3017_), .B(_3025_), .Q(_3026_) );
NA2X1 NA2X1_864 ( .gnd!(gnd!), .vdd!(vdd!), .A(_3024_), .B(_3022_), .Q(_3027_) );
NA2I1X1 NA2I1X1_126 ( .gnd!(gnd!), .vdd!(vdd!), .AN(_3017_), .B(_3027_), .Q(_3028_) );
AND2X2 AND2X2_90 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_IDEC1_cu_jalr_inst_bF_buf2), .B(ALU_r_19_), .Q(_3029_) );
AN31X1 AN31X1_86 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2686__bF_buf1), .B(_3026_), .C(_3028_), .D(_3029_), .Q(_3030_) );
MU2IX1 MU2IX1_120 ( .gnd!(gnd!), .vdd!(vdd!), .IN0(_3030_), .IN1(_3016_), .Q(_3031_), .S(_2647__bF_buf4) );
MU2X1 MU2X1_246 ( .gnd!(gnd!), .vdd!(vdd!), .IN0(_3031_), .IN1(PCU_ePC_19_), .Q(_2642__19_), .S(_2643__bF_buf3) );
NA2X1 NA2X1_865 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2643__bF_buf0), .B(PCU_ePC_20_), .Q(_3032_) );
AND2X2 AND2X2_91 ( .gnd!(gnd!), .vdd!(vdd!), .A(_3007_), .B(_3010_), .Q(_3033_) );
NO2X1 NO2X1_365 ( .gnd!(gnd!), .vdd!(vdd!), .A(_3019_), .B(_3021_), .Q(_3034_) );
ON21X1 ON21X1_356 ( .gnd!(gnd!), .vdd!(vdd!), .A(_3034_), .B(_3010_), .C(_3022_), .Q(_3035_) );
AN31X1 AN31X1_87 ( .gnd!(gnd!), .vdd!(vdd!), .A(_3003_), .B(_3025_), .C(_3033_), .D(_3035_), .Q(_3036_) );
NO2X1 NO2X1_366 ( .gnd!(gnd!), .vdd!(vdd!), .A(_3011_), .B(_3027_), .Q(_3037_) );
NA2X1 NA2X1_866 ( .gnd!(gnd!), .vdd!(vdd!), .A(_3001_), .B(_3037_), .Q(_3038_) );
ON21X1 ON21X1_357 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2981_), .B(_3038_), .C(_3036_), .Q(_3039_) );
INX1 INX1_224 ( .gnd!(gnd!), .vdd!(vdd!), .A(PC_20_), .Q(_3040_) );
NA2X1 NA2X1_867 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_cu_pc_s2_bF_buf7), .B(I1_20_), .Q(_3041_) );
NO2X1 NO2X1_367 ( .gnd!(gnd!), .vdd!(vdd!), .A(PC1_20_), .B(_2650__bF_buf0), .Q(_3042_) );
AO211X4 AO211X4_3 ( .gnd!(gnd!), .vdd!(vdd!), .A(_3040_), .B(_2650__bF_buf0), .C(_3041_), .D(_3042_), .Q(_3043_) );
MU2IX1 MU2IX1_121 ( .gnd!(gnd!), .vdd!(vdd!), .IN0(PC1_20_), .IN1(PC_20_), .Q(_3044_), .S(_2650__bF_buf0) );
NA2X1 NA2X1_868 ( .gnd!(gnd!), .vdd!(vdd!), .A(_3044_), .B(_3041_), .Q(_3045_) );
NA2X1 NA2X1_869 ( .gnd!(gnd!), .vdd!(vdd!), .A(_3045_), .B(_3043_), .Q(_3046_) );
EN2X1 EN2X1_28 ( .gnd!(gnd!), .vdd!(vdd!), .A(_3039_), .B(_3046_), .Q(_3047_) );
MU2X1 MU2X1_247 ( .gnd!(gnd!), .vdd!(vdd!), .IN0(_3047_), .IN1(ALU_r_20_), .Q(_3048_), .S(CTRL_IDEC1_cu_jalr_inst_bF_buf1) );
NO2X1 NO2X1_368 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2647__bF_buf4), .B(_3048_), .Q(_3049_) );
NO2X1 NO2X1_369 ( .gnd!(gnd!), .vdd!(vdd!), .A(PC_20_), .B(_2646__bF_buf1), .Q(_3050_) );
ON31X1 ON31X1_94 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2643__bF_buf0), .B(_3050_), .C(_3049_), .D(_3032_), .Q(_2642__20_) );
NA2X1 NA2X1_870 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_IDEC1_cu_jalr_inst_bF_buf2), .B(ALU_r_21_), .Q(_3051_) );
NO2X1 NO2X1_370 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2963_), .B(_2966_), .Q(_3052_) );
NO2X1 NO2X1_371 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2986_), .B(_2990_), .Q(_3053_) );
AN21X1 AN21X1_181 ( .gnd!(gnd!), .vdd!(vdd!), .A(_3052_), .B(_2991_), .C(_3053_), .Q(_3054_) );
NA2I1X1 NA2I1X1_127 ( .gnd!(gnd!), .vdd!(vdd!), .AN(_3010_), .B(_3024_), .Q(_3055_) );
ON311X1 ON311X1_17 ( .gnd!(gnd!), .vdd!(vdd!), .A(_3011_), .B(_3034_), .C(_3054_), .D(_3022_), .E(_3055_), .Q(_3056_) );
AN31X1 AN31X1_88 ( .gnd!(gnd!), .vdd!(vdd!), .A(_3001_), .B(_3037_), .C(_2961_), .D(_3056_), .Q(_3057_) );
NA2X1 NA2X1_871 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_cu_pc_s2_bF_buf7), .B(I1_21_), .Q(_3058_) );
INX1 INX1_225 ( .gnd!(gnd!), .vdd!(vdd!), .A(_3058_), .Q(_3059_) );
MU2IX1 MU2IX1_122 ( .gnd!(gnd!), .vdd!(vdd!), .IN0(PC1_21_), .IN1(PC_21_), .Q(_3060_), .S(_2650__bF_buf0) );
NO2X1 NO2X1_372 ( .gnd!(gnd!), .vdd!(vdd!), .A(_3059_), .B(_3060_), .Q(_3061_) );
INX1 INX1_226 ( .gnd!(gnd!), .vdd!(vdd!), .A(PC_21_), .Q(_3062_) );
NO2X1 NO2X1_373 ( .gnd!(gnd!), .vdd!(vdd!), .A(PC1_21_), .B(_2650__bF_buf0), .Q(_3063_) );
AN21X1 AN21X1_182 ( .gnd!(gnd!), .vdd!(vdd!), .A(_3062_), .B(_2650__bF_buf0), .C(_3063_), .Q(_3064_) );
NO2X1 NO2X1_374 ( .gnd!(gnd!), .vdd!(vdd!), .A(_3058_), .B(_3064_), .Q(_3065_) );
ON211X1 ON211X1_124 ( .gnd!(gnd!), .vdd!(vdd!), .A(_3061_), .B(_3065_), .C(_3043_), .D(_3045_), .Q(_3066_) );
NO2X1 NO2X1_375 ( .gnd!(gnd!), .vdd!(vdd!), .A(_3066_), .B(_3057_), .Q(_3067_) );
NO2X1 NO2X1_376 ( .gnd!(gnd!), .vdd!(vdd!), .A(_3041_), .B(_3044_), .Q(_3068_) );
NA2X1 NA2X1_872 ( .gnd!(gnd!), .vdd!(vdd!), .A(_3064_), .B(_3059_), .Q(_3069_) );
NA2X1 NA2X1_873 ( .gnd!(gnd!), .vdd!(vdd!), .A(_3060_), .B(_3058_), .Q(_3070_) );
AN221X1 AN221X1_9 ( .gnd!(gnd!), .vdd!(vdd!), .A(_3069_), .B(_3070_), .C(_3039_), .D(_3045_), .E(_3068_), .Q(_3071_) );
NO2X1 NO2X1_377 ( .gnd!(gnd!), .vdd!(vdd!), .A(_3058_), .B(_3060_), .Q(_3072_) );
NO2X1 NO2X1_378 ( .gnd!(gnd!), .vdd!(vdd!), .A(_3059_), .B(_3064_), .Q(_3073_) );
ON31X1 ON31X1_95 ( .gnd!(gnd!), .vdd!(vdd!), .A(_3043_), .B(_3073_), .C(_3072_), .D(_2686__bF_buf1), .Q(_3074_) );
ON31X1 ON31X1_96 ( .gnd!(gnd!), .vdd!(vdd!), .A(_3067_), .B(_3074_), .C(_3071_), .D(_3051_), .Q(_3075_) );
MU2X1 MU2X1_248 ( .gnd!(gnd!), .vdd!(vdd!), .IN0(_3075_), .IN1(PC_21_), .Q(_3076_), .S(_2647__bF_buf4) );
MU2X1 MU2X1_249 ( .gnd!(gnd!), .vdd!(vdd!), .IN0(_3076_), .IN1(PCU_ePC_21_), .Q(_2642__21_), .S(_2643__bF_buf3) );
NA2X1 NA2X1_874 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2643__bF_buf0), .B(PCU_ePC_22_), .Q(_3077_) );
AND2X2 AND2X2_92 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_IDEC1_cu_jalr_inst_bF_buf0), .B(ALU_r_22_), .Q(_3078_) );
AN21X1 AN21X1_183 ( .gnd!(gnd!), .vdd!(vdd!), .A(_3068_), .B(_3070_), .C(_3072_), .Q(_3079_) );
ON21X1 ON21X1_358 ( .gnd!(gnd!), .vdd!(vdd!), .A(_3057_), .B(_3066_), .C(_3079_), .Q(_3080_) );
NA2X1 NA2X1_875 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_cu_pc_s2_bF_buf4), .B(I1_22_), .Q(_3081_) );
MU2X1 MU2X1_250 ( .gnd!(gnd!), .vdd!(vdd!), .IN0(PC1_22_), .IN1(PC_22_), .Q(_3082_), .S(_2650__bF_buf5) );
NA2X1 NA2X1_876 ( .gnd!(gnd!), .vdd!(vdd!), .A(_3082_), .B(_3081_), .Q(_3083_) );
INX1 INX1_227 ( .gnd!(gnd!), .vdd!(vdd!), .A(_3081_), .Q(_3084_) );
MU2IX1 MU2IX1_123 ( .gnd!(gnd!), .vdd!(vdd!), .IN0(PC1_22_), .IN1(PC_22_), .Q(_3085_), .S(_2650__bF_buf5) );
NA2X1 NA2X1_877 ( .gnd!(gnd!), .vdd!(vdd!), .A(_3085_), .B(_3084_), .Q(_3086_) );
AND2X2 AND2X2_93 ( .gnd!(gnd!), .vdd!(vdd!), .A(_3083_), .B(_3086_), .Q(_3087_) );
NA2I1X1 NA2I1X1_128 ( .gnd!(gnd!), .vdd!(vdd!), .AN(_3080_), .B(_3087_), .Q(_3088_) );
INX1 INX1_228 ( .gnd!(gnd!), .vdd!(vdd!), .A(_3087_), .Q(_3089_) );
NA2X1 NA2X1_878 ( .gnd!(gnd!), .vdd!(vdd!), .A(_3080_), .B(_3089_), .Q(_3090_) );
AND3X4 AND3X4_17 ( .gnd!(gnd!), .vdd!(vdd!), .A(_3088_), .B(_2686__bF_buf1), .C(_3090_), .Q(_3091_) );
NO3X1 NO3X1_22 ( .gnd!(gnd!), .vdd!(vdd!), .A(_3091_), .B(_2647__bF_buf0), .C(_3078_), .Q(_3092_) );
NO2X1 NO2X1_379 ( .gnd!(gnd!), .vdd!(vdd!), .A(PC_22_), .B(_2646__bF_buf1), .Q(_3093_) );
ON31X1 ON31X1_97 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2643__bF_buf0), .B(_3093_), .C(_3092_), .D(_3077_), .Q(_2642__22_) );
NA2X1 NA2X1_879 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2643__bF_buf3), .B(PCU_ePC_23_), .Q(_3094_) );
NA2I1X1 NA2I1X1_129 ( .gnd!(gnd!), .vdd!(vdd!), .AN(ALU_r_23_), .B(CTRL_IDEC1_cu_jalr_inst_bF_buf1), .Q(_3095_) );
NA2X1 NA2X1_880 ( .gnd!(gnd!), .vdd!(vdd!), .A(_3082_), .B(_3084_), .Q(_3096_) );
INX1 INX1_229 ( .gnd!(gnd!), .vdd!(vdd!), .A(PC_23_), .Q(_3097_) );
NA2X1 NA2X1_881 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_cu_pc_s2_bF_buf4), .B(I1_23_), .Q(_3098_) );
NO2X1 NO2X1_380 ( .gnd!(gnd!), .vdd!(vdd!), .A(PC1_23_), .B(_2650__bF_buf7), .Q(_3099_) );
AO211X4 AO211X4_4 ( .gnd!(gnd!), .vdd!(vdd!), .A(_3097_), .B(_2650__bF_buf5), .C(_3098_), .D(_3099_), .Q(_3100_) );
MU2IX1 MU2IX1_124 ( .gnd!(gnd!), .vdd!(vdd!), .IN0(PC1_23_), .IN1(PC_23_), .Q(_3101_), .S(_2650__bF_buf5) );
NA2X1 NA2X1_882 ( .gnd!(gnd!), .vdd!(vdd!), .A(_3101_), .B(_3098_), .Q(_3102_) );
NA2X1 NA2X1_883 ( .gnd!(gnd!), .vdd!(vdd!), .A(_3102_), .B(_3100_), .Q(_3103_) );
AN21X1 AN21X1_184 ( .gnd!(gnd!), .vdd!(vdd!), .A(_3090_), .B(_3096_), .C(_3103_), .Q(_3104_) );
NO2X1 NO2X1_381 ( .gnd!(gnd!), .vdd!(vdd!), .A(_3081_), .B(_3085_), .Q(_3105_) );
AN221X1 AN221X1_10 ( .gnd!(gnd!), .vdd!(vdd!), .A(_3100_), .B(_3102_), .C(_3080_), .D(_3089_), .E(_3105_), .Q(_3106_) );
ON21X1 ON21X1_359 ( .gnd!(gnd!), .vdd!(vdd!), .A(_3104_), .B(_3106_), .C(_2686__bF_buf1), .Q(_3107_) );
NO2X1 NO2X1_382 ( .gnd!(gnd!), .vdd!(vdd!), .A(_3097_), .B(_2646__bF_buf3), .Q(_3108_) );
AN31X1 AN31X1_89 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2646__bF_buf3), .B(_3095_), .C(_3107_), .D(_3108_), .Q(_3109_) );
ON21X1 ON21X1_360 ( .gnd!(gnd!), .vdd!(vdd!), .A(_3109_), .B(_2643__bF_buf3), .C(_3094_), .Q(_2642__23_) );
NO3X1 NO3X1_23 ( .gnd!(gnd!), .vdd!(vdd!), .A(_3087_), .B(_3066_), .C(_3103_), .Q(_3110_) );
NO2X1 NO2X1_383 ( .gnd!(gnd!), .vdd!(vdd!), .A(_3098_), .B(_3101_), .Q(_3111_) );
AN21X1 AN21X1_185 ( .gnd!(gnd!), .vdd!(vdd!), .A(_3105_), .B(_3102_), .C(_3111_), .Q(_3112_) );
ON31X1 ON31X1_98 ( .gnd!(gnd!), .vdd!(vdd!), .A(_3103_), .B(_3079_), .C(_3087_), .D(_3112_), .Q(_3113_) );
AN21X1 AN21X1_186 ( .gnd!(gnd!), .vdd!(vdd!), .A(_3110_), .B(_3056_), .C(_3113_), .Q(_3114_) );
NA2I1X1 NA2I1X1_130 ( .gnd!(gnd!), .vdd!(vdd!), .AN(_3038_), .B(_3110_), .Q(_3115_) );
ON21X1 ON21X1_361 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2981_), .B(_3115_), .C(_3114_), .Q(_3116_) );
AND2X2 AND2X2_94 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_cu_pc_s2_bF_buf2), .B(I1_24_), .Q(_3118_) );
MU2X1 MU2X1_251 ( .gnd!(gnd!), .vdd!(vdd!), .IN0(PC1_24_), .IN1(PC_24_), .Q(_3119_), .S(_2650__bF_buf6) );
OR2X2 OR2X2_25 ( .gnd!(gnd!), .vdd!(vdd!), .A(_3119_), .B(_3118_), .Q(_3120_) );
NA2X1 NA2X1_884 ( .gnd!(gnd!), .vdd!(vdd!), .A(_3119_), .B(_3118_), .Q(_3121_) );
NA2X1 NA2X1_885 ( .gnd!(gnd!), .vdd!(vdd!), .A(_3120_), .B(_3121_), .Q(_3122_) );
INX1 INX1_230 ( .gnd!(gnd!), .vdd!(vdd!), .A(_3122_), .Q(_3123_) );
NO2X1 NO2X1_384 ( .gnd!(gnd!), .vdd!(vdd!), .A(_3123_), .B(_3116_), .Q(_3124_) );
AN21X1 AN21X1_187 ( .gnd!(gnd!), .vdd!(vdd!), .A(_3083_), .B(_3086_), .C(_3103_), .Q(_3125_) );
NA2I1X1 NA2I1X1_131 ( .gnd!(gnd!), .vdd!(vdd!), .AN(_3066_), .B(_3125_), .Q(_3126_) );
ON21X1 ON21X1_362 ( .gnd!(gnd!), .vdd!(vdd!), .A(_3073_), .B(_3043_), .C(_3069_), .Q(_3127_) );
ON21X1 ON21X1_363 ( .gnd!(gnd!), .vdd!(vdd!), .A(_3103_), .B(_3096_), .C(_3100_), .Q(_3128_) );
AN21X1 AN21X1_188 ( .gnd!(gnd!), .vdd!(vdd!), .A(_3125_), .B(_3127_), .C(_3128_), .Q(_3129_) );
ON21X1 ON21X1_364 ( .gnd!(gnd!), .vdd!(vdd!), .A(_3036_), .B(_3126_), .C(_3129_), .Q(_3130_) );
NO2X1 NO2X1_385 ( .gnd!(gnd!), .vdd!(vdd!), .A(_3038_), .B(_3126_), .Q(_3131_) );
AN21X1 AN21X1_189 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2961_), .B(_3131_), .C(_3130_), .Q(_3132_) );
NO2X1 NO2X1_386 ( .gnd!(gnd!), .vdd!(vdd!), .A(_3122_), .B(_3132_), .Q(_3133_) );
NA2X1 NA2X1_886 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_IDEC1_cu_jalr_inst_bF_buf3), .B(ALU_r_24_), .Q(_3134_) );
ON31X1 ON31X1_99 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_IDEC1_cu_jalr_inst_bF_buf0), .B(_3133_), .C(_3124_), .D(_3134_), .Q(_3135_) );
MU2X1 MU2X1_252 ( .gnd!(gnd!), .vdd!(vdd!), .IN0(_3135_), .IN1(PC_24_), .Q(_3136_), .S(_2647__bF_buf2) );
MU2X1 MU2X1_253 ( .gnd!(gnd!), .vdd!(vdd!), .IN0(_3136_), .IN1(PCU_ePC_24_), .Q(_2642__24_), .S(_2643__bF_buf5) );
NA2X1 NA2X1_887 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_IDEC1_cu_jalr_inst_bF_buf3), .B(ALU_r_25_), .Q(_3137_) );
NA2X1 NA2X1_888 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_cu_pc_s2_bF_buf2), .B(I1_25_), .Q(_3138_) );
MU2X1 MU2X1_254 ( .gnd!(gnd!), .vdd!(vdd!), .IN0(PC1_25_), .IN1(PC_25_), .Q(_3139_), .S(_2650__bF_buf6) );
NA2I1X1 NA2I1X1_132 ( .gnd!(gnd!), .vdd!(vdd!), .AN(_3138_), .B(_3139_), .Q(_3140_) );
MU2IX1 MU2IX1_125 ( .gnd!(gnd!), .vdd!(vdd!), .IN0(PC1_25_), .IN1(PC_25_), .Q(_3141_), .S(_2650__bF_buf6) );
NA2X1 NA2X1_889 ( .gnd!(gnd!), .vdd!(vdd!), .A(_3141_), .B(_3138_), .Q(_3142_) );
NA2X1 NA2X1_890 ( .gnd!(gnd!), .vdd!(vdd!), .A(_3140_), .B(_3142_), .Q(_3143_) );
NO2X1 NO2X1_387 ( .gnd!(gnd!), .vdd!(vdd!), .A(_3121_), .B(_3143_), .Q(_3144_) );
NO2X1 NO2X1_388 ( .gnd!(gnd!), .vdd!(vdd!), .A(_3143_), .B(_3122_), .Q(_3145_) );
INX1 INX1_231 ( .gnd!(gnd!), .vdd!(vdd!), .A(_3145_), .Q(_3146_) );
NA2X1 NA2X1_891 ( .gnd!(gnd!), .vdd!(vdd!), .A(_3143_), .B(_3121_), .Q(_3147_) );
ON22X1 ON22X1_84 ( .gnd!(gnd!), .vdd!(vdd!), .A(_3133_), .B(_3147_), .C(_3132_), .D(_3146_), .Q(_3148_) );
ON31X1 ON31X1_100 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_IDEC1_cu_jalr_inst_bF_buf0), .B(_3144_), .C(_3148_), .D(_3137_), .Q(_3149_) );
MU2X1 MU2X1_255 ( .gnd!(gnd!), .vdd!(vdd!), .IN0(_3149_), .IN1(PC_25_), .Q(_3150_), .S(_2647__bF_buf3) );
MU2X1 MU2X1_256 ( .gnd!(gnd!), .vdd!(vdd!), .IN0(_3150_), .IN1(PCU_ePC_25_), .Q(_2642__25_), .S(_2643__bF_buf4) );
NA2X1 NA2X1_892 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2643__bF_buf5), .B(PCU_ePC_26_), .Q(_3151_) );
AND2X2 AND2X2_95 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_IDEC1_cu_jalr_inst_bF_buf3), .B(ALU_r_26_), .Q(_3152_) );
NO2I1X1 NO2I1X1_56 ( .gnd!(gnd!), .vdd!(vdd!), .AN(_3140_), .B(_3144_), .Q(_3153_) );
ON21X1 ON21X1_365 ( .gnd!(gnd!), .vdd!(vdd!), .A(_3132_), .B(_3146_), .C(_3153_), .Q(_3154_) );
AND2X2 AND2X2_96 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_cu_pc_s2_bF_buf2), .B(I1_26_), .Q(_3155_) );
MU2IX1 MU2IX1_126 ( .gnd!(gnd!), .vdd!(vdd!), .IN0(PC1_26_), .IN1(PC_26_), .Q(_3156_), .S(_2650__bF_buf1) );
NA2I1X1 NA2I1X1_133 ( .gnd!(gnd!), .vdd!(vdd!), .AN(_3155_), .B(_3156_), .Q(_3157_) );
NA2I1X1 NA2I1X1_134 ( .gnd!(gnd!), .vdd!(vdd!), .AN(_3156_), .B(_3155_), .Q(_3158_) );
AND2X2 AND2X2_97 ( .gnd!(gnd!), .vdd!(vdd!), .A(_3158_), .B(_3157_), .Q(_3159_) );
NA2X1 NA2X1_893 ( .gnd!(gnd!), .vdd!(vdd!), .A(_3154_), .B(_3159_), .Q(_3160_) );
OR2X2 OR2X2_26 ( .gnd!(gnd!), .vdd!(vdd!), .A(_3154_), .B(_3159_), .Q(_3161_) );
AND3X4 AND3X4_18 ( .gnd!(gnd!), .vdd!(vdd!), .A(_3161_), .B(_2686__bF_buf2), .C(_3160_), .Q(_3162_) );
NO3X1 NO3X1_24 ( .gnd!(gnd!), .vdd!(vdd!), .A(_3162_), .B(_2647__bF_buf3), .C(_3152_), .Q(_3163_) );
NO2X1 NO2X1_389 ( .gnd!(gnd!), .vdd!(vdd!), .A(PC_26_), .B(_2646__bF_buf1), .Q(_3164_) );
ON31X1 ON31X1_101 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2643__bF_buf4), .B(_3164_), .C(_3163_), .D(_3151_), .Q(_2642__26_) );
NA2X1 NA2X1_894 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2643__bF_buf4), .B(PCU_ePC_27_), .Q(_3165_) );
NA2I1X1 NA2I1X1_135 ( .gnd!(gnd!), .vdd!(vdd!), .AN(ALU_r_27_), .B(CTRL_IDEC1_cu_jalr_inst_bF_buf0), .Q(_3166_) );
AND2X2 AND2X2_98 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_cu_pc_s2_bF_buf2), .B(I1_27_), .Q(_3167_) );
MU2IX1 MU2IX1_127 ( .gnd!(gnd!), .vdd!(vdd!), .IN0(PC1_27_), .IN1(PC_27_), .Q(_3168_), .S(_2650__bF_buf6) );
NA2I1X1 NA2I1X1_136 ( .gnd!(gnd!), .vdd!(vdd!), .AN(_3168_), .B(_3167_), .Q(_3169_) );
NA2I1X1 NA2I1X1_137 ( .gnd!(gnd!), .vdd!(vdd!), .AN(_3167_), .B(_3168_), .Q(_3170_) );
NA2X1 NA2X1_895 ( .gnd!(gnd!), .vdd!(vdd!), .A(_3169_), .B(_3170_), .Q(_3171_) );
AN21X1 AN21X1_190 ( .gnd!(gnd!), .vdd!(vdd!), .A(_3160_), .B(_3158_), .C(_3171_), .Q(_3172_) );
AND3X4 AND3X4_19 ( .gnd!(gnd!), .vdd!(vdd!), .A(_3160_), .B(_3158_), .C(_3171_), .Q(_3173_) );
ON21X1 ON21X1_366 ( .gnd!(gnd!), .vdd!(vdd!), .A(_3173_), .B(_3172_), .C(_2686__bF_buf2), .Q(_3174_) );
INX1 INX1_232 ( .gnd!(gnd!), .vdd!(vdd!), .A(PC_27_), .Q(_3175_) );
NO2X1 NO2X1_390 ( .gnd!(gnd!), .vdd!(vdd!), .A(_3175_), .B(_2646__bF_buf0), .Q(_3176_) );
AN31X1 AN31X1_90 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2646__bF_buf0), .B(_3166_), .C(_3174_), .D(_3176_), .Q(_3177_) );
ON21X1 ON21X1_367 ( .gnd!(gnd!), .vdd!(vdd!), .A(_3177_), .B(_2643__bF_buf2), .C(_3165_), .Q(_2642__27_) );
NA2X1 NA2X1_896 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2643__bF_buf2), .B(PCU_ePC_28_), .Q(_3178_) );
NA2I1X1 NA2I1X1_138 ( .gnd!(gnd!), .vdd!(vdd!), .AN(_3171_), .B(_3159_), .Q(_3179_) );
NO2X1 NO2X1_391 ( .gnd!(gnd!), .vdd!(vdd!), .A(_3179_), .B(_3146_), .Q(_3180_) );
ON221X1 ON221X1_21 ( .gnd!(gnd!), .vdd!(vdd!), .A(_3158_), .B(_3171_), .C(_3153_), .D(_3179_), .E(_3169_), .Q(_3181_) );
AN21X1 AN21X1_191 ( .gnd!(gnd!), .vdd!(vdd!), .A(_3116_), .B(_3180_), .C(_3181_), .Q(_3182_) );
NA2X1 NA2X1_897 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_cu_pc_s2_bF_buf2), .B(I1_28_), .Q(_3183_) );
MU2IX1 MU2IX1_128 ( .gnd!(gnd!), .vdd!(vdd!), .IN0(PC1_28_), .IN1(PC_28_), .Q(_3184_), .S(_2650__bF_buf6) );
NO2X1 NO2X1_392 ( .gnd!(gnd!), .vdd!(vdd!), .A(_3183_), .B(_3184_), .Q(_3185_) );
INX1 INX1_233 ( .gnd!(gnd!), .vdd!(vdd!), .A(_3185_), .Q(_3186_) );
NA2X1 NA2X1_898 ( .gnd!(gnd!), .vdd!(vdd!), .A(_3184_), .B(_3183_), .Q(_3187_) );
NA2X1 NA2X1_899 ( .gnd!(gnd!), .vdd!(vdd!), .A(_3186_), .B(_3187_), .Q(_3188_) );
NO2X1 NO2X1_393 ( .gnd!(gnd!), .vdd!(vdd!), .A(_3188_), .B(_3182_), .Q(_3189_) );
NA2I1X1 NA2I1X1_139 ( .gnd!(gnd!), .vdd!(vdd!), .AN(_3179_), .B(_3145_), .Q(_3190_) );
OA221X1 OA221X1_2 ( .gnd!(gnd!), .vdd!(vdd!), .A(_3158_), .B(_3171_), .C(_3153_), .D(_3179_), .E(_3169_), .Q(_3191_) );
ON21X1 ON21X1_368 ( .gnd!(gnd!), .vdd!(vdd!), .A(_3132_), .B(_3190_), .C(_3191_), .Q(_3192_) );
INX1 INX1_234 ( .gnd!(gnd!), .vdd!(vdd!), .A(_3188_), .Q(_3193_) );
NO2X1 NO2X1_394 ( .gnd!(gnd!), .vdd!(vdd!), .A(_3193_), .B(_3192_), .Q(_3194_) );
NA2X1 NA2X1_900 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_IDEC1_cu_jalr_inst_bF_buf5), .B(ALU_r_28_), .Q(_3195_) );
ON31X1 ON31X1_102 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_IDEC1_cu_jalr_inst_bF_buf3), .B(_3194_), .C(_3189_), .D(_3195_), .Q(_3196_) );
NO2X1 NO2X1_395 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2647__bF_buf3), .B(_3196_), .Q(_3197_) );
NO2X1 NO2X1_396 ( .gnd!(gnd!), .vdd!(vdd!), .A(PC_28_), .B(_2646__bF_buf0), .Q(_3198_) );
ON31X1 ON31X1_103 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2643__bF_buf2), .B(_3198_), .C(_3197_), .D(_3178_), .Q(_2642__28_) );
NA2X1 NA2X1_901 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2643__bF_buf1), .B(PCU_ePC_29_), .Q(_3199_) );
NA2X1 NA2X1_902 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_IDEC1_cu_jalr_inst_bF_buf5), .B(ALU_r_29_), .Q(_3200_) );
AND2X2 AND2X2_99 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_cu_pc_s2_bF_buf1), .B(I1_29_), .Q(_3201_) );
MU2X1 MU2X1_257 ( .gnd!(gnd!), .vdd!(vdd!), .IN0(PC1_29_), .IN1(PC_29_), .Q(_3202_), .S(_2650__bF_buf2) );
AND2X2 AND2X2_100 ( .gnd!(gnd!), .vdd!(vdd!), .A(_3202_), .B(_3201_), .Q(_3203_) );
NO2X1 NO2X1_397 ( .gnd!(gnd!), .vdd!(vdd!), .A(_3201_), .B(_3202_), .Q(_3204_) );
NO2X1 NO2X1_398 ( .gnd!(gnd!), .vdd!(vdd!), .A(_3204_), .B(_3203_), .Q(_3205_) );
NA2X1 NA2X1_903 ( .gnd!(gnd!), .vdd!(vdd!), .A(_3205_), .B(_3185_), .Q(_3206_) );
NA2X1 NA2X1_904 ( .gnd!(gnd!), .vdd!(vdd!), .A(_3206_), .B(_2686__bF_buf3), .Q(_3207_) );
NA2X1 NA2X1_905 ( .gnd!(gnd!), .vdd!(vdd!), .A(_3193_), .B(_3205_), .Q(_3208_) );
ON32X1 ON32X1_7 ( .gnd!(gnd!), .vdd!(vdd!), .A(_3185_), .B(_3205_), .C(_3189_), .D(_3182_), .E(_3208_), .Q(_3209_) );
ON21X1 ON21X1_369 ( .gnd!(gnd!), .vdd!(vdd!), .A(_3209_), .B(_3207_), .C(_3200_), .Q(_3210_) );
INX1 INX1_235 ( .gnd!(gnd!), .vdd!(vdd!), .A(PC_29_), .Q(_3211_) );
NA2X1 NA2X1_906 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2647__bF_buf1), .B(_3211_), .Q(_3212_) );
ON211X1 ON211X1_125 ( .gnd!(gnd!), .vdd!(vdd!), .A(_3210_), .B(_2647__bF_buf1), .C(CTRL_cu_ld_epc), .D(_3212_), .Q(_3213_) );
NA2X1 NA2X1_907 ( .gnd!(gnd!), .vdd!(vdd!), .A(_3213_), .B(_3199_), .Q(_2642__29_) );
INX1 INX1_236 ( .gnd!(gnd!), .vdd!(vdd!), .A(_3208_), .Q(_3214_) );
NA2I1X1 NA2I1X1_140 ( .gnd!(gnd!), .vdd!(vdd!), .AN(_3203_), .B(_3206_), .Q(_3215_) );
AN21X1 AN21X1_192 ( .gnd!(gnd!), .vdd!(vdd!), .A(_3192_), .B(_3214_), .C(_3215_), .Q(_3216_) );
NA2X1 NA2X1_908 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_cu_pc_s2_bF_buf1), .B(I1_30_), .Q(_3217_) );
INX1 INX1_237 ( .gnd!(gnd!), .vdd!(vdd!), .A(_3217_), .Q(_3218_) );
MU2X1 MU2X1_258 ( .gnd!(gnd!), .vdd!(vdd!), .IN0(PC1_30_), .IN1(PC_30_), .Q(_3219_), .S(_2650__bF_buf6) );
NO2X1 NO2X1_399 ( .gnd!(gnd!), .vdd!(vdd!), .A(_3218_), .B(_3219_), .Q(_3220_) );
NA2X1 NA2X1_909 ( .gnd!(gnd!), .vdd!(vdd!), .A(_3219_), .B(_3218_), .Q(_3221_) );
NA2I1X1 NA2I1X1_141 ( .gnd!(gnd!), .vdd!(vdd!), .AN(_3220_), .B(_3221_), .Q(_3222_) );
NA2X1 NA2X1_910 ( .gnd!(gnd!), .vdd!(vdd!), .A(_3216_), .B(_3222_), .Q(_3223_) );
INX1 INX1_238 ( .gnd!(gnd!), .vdd!(vdd!), .A(_3215_), .Q(_3224_) );
ON21X1 ON21X1_370 ( .gnd!(gnd!), .vdd!(vdd!), .A(_3182_), .B(_3208_), .C(_3224_), .Q(_3225_) );
INX1 INX1_239 ( .gnd!(gnd!), .vdd!(vdd!), .A(_3222_), .Q(_3226_) );
NA2X1 NA2X1_911 ( .gnd!(gnd!), .vdd!(vdd!), .A(_3225_), .B(_3226_), .Q(_3227_) );
NA2X1 NA2X1_912 ( .gnd!(gnd!), .vdd!(vdd!), .A(_3227_), .B(_3223_), .Q(_3228_) );
NA2X1 NA2X1_913 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_IDEC1_cu_jalr_inst_bF_buf4), .B(ALU_r_30_), .Q(_3229_) );
ON211X1 ON211X1_126 ( .gnd!(gnd!), .vdd!(vdd!), .A(_3228_), .B(CTRL_IDEC1_cu_jalr_inst_bF_buf0), .C(_2646__bF_buf2), .D(_3229_), .Q(_3230_) );
NO2X1 NO2X1_400 ( .gnd!(gnd!), .vdd!(vdd!), .A(PC_30_), .B(_2646__bF_buf2), .Q(_3231_) );
NO2X1 NO2X1_401 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2643__bF_buf2), .B(_3231_), .Q(_3232_) );
AO22X2 AO22X2_42 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2643__bF_buf2), .B(PCU_ePC_30_), .C(_3230_), .D(_3232_), .Q(_2642__30_) );
NA2X1 NA2X1_914 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2643__bF_buf2), .B(PCU_ePC_31_), .Q(_3233_) );
ON21X1 ON21X1_371 ( .gnd!(gnd!), .vdd!(vdd!), .A(_3216_), .B(_3220_), .C(_3221_), .Q(_3234_) );
AND2X2 AND2X2_101 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_cu_pc_s2_bF_buf1), .B(I1_31_), .Q(_3235_) );
MU2IX1 MU2IX1_129 ( .gnd!(gnd!), .vdd!(vdd!), .IN0(PC1_31_), .IN1(PC_31_), .Q(_3236_), .S(_2650__bF_buf6) );
EN2X1 EN2X1_29 ( .gnd!(gnd!), .vdd!(vdd!), .A(_3236_), .B(_3235_), .Q(_3237_) );
NA2X1 NA2X1_915 ( .gnd!(gnd!), .vdd!(vdd!), .A(_3234_), .B(_3237_), .Q(_3238_) );
NA3I1X1 NA3I1X1_129 ( .gnd!(gnd!), .vdd!(vdd!), .AN(_3237_), .B(_3221_), .C(_3227_), .Q(_3239_) );
INX1 INX1_240 ( .gnd!(gnd!), .vdd!(vdd!), .A(ALU_r_31_), .Q(_3240_) );
NO2X1 NO2X1_402 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2686__bF_buf3), .B(_3240_), .Q(_3241_) );
AN311X1 AN311X1_4 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2686__bF_buf3), .B(_3239_), .C(_3238_), .D(_2647__bF_buf3), .E(_3241_), .Q(_3242_) );
ON21X1 ON21X1_372 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2646__bF_buf2), .B(PC_31_), .C(CTRL_cu_ld_epc), .Q(_3243_) );
ON21X1 ON21X1_373 ( .gnd!(gnd!), .vdd!(vdd!), .A(_3242_), .B(_3243_), .C(_3233_), .Q(_2642__31_) );
NO2X1 NO2X1_403 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_cu_pc_s4_bF_buf2), .B(CTRL_cu_pc_s0), .Q(_3244_) );
AO22X2 AO22X2_43 ( .gnd!(gnd!), .vdd!(vdd!), .A(PCU_ePC_0_), .B(CTRL_cu_pc_s4_bF_buf3), .C(_2657_), .D(_3244__bF_buf1), .Q(_3245_) );
NA2I1X2 NA2I1X2_4 ( .gnd!(gnd!), .vdd!(vdd!), .AN(CTRL_cu_ext_hold_bF_buf4), .B(CTRL_cyc_bF_buf0_bF_buf0), .Q(_3246_) );
MU2X1 MU2X1_259 ( .gnd!(gnd!), .vdd!(vdd!), .IN0(_3245_), .IN1(PC_0_), .Q(_2641__0_), .S(_3246__bF_buf1) );
INX2 INX2_15 ( .gnd!(gnd!), .vdd!(vdd!), .A(_3246__bF_buf2), .Q(_3247_) );
NO2X1 NO2X1_404 ( .gnd!(gnd!), .vdd!(vdd!), .A(PC_1_), .B(_3247__bF_buf3), .Q(_3248_) );
NA2X1 NA2X1_916 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2668_), .B(_3244__bF_buf4), .Q(_3249_) );
NA2X1 NA2X1_917 ( .gnd!(gnd!), .vdd!(vdd!), .A(PCU_ePC_1_), .B(CTRL_cu_pc_s4_bF_buf1), .Q(_3250_) );
AN31X1 AN31X1_91 ( .gnd!(gnd!), .vdd!(vdd!), .A(_3247__bF_buf3), .B(_3250_), .C(_3249_), .D(_3248_), .Q(_2641__1_) );
NO2X1 NO2X1_405 ( .gnd!(gnd!), .vdd!(vdd!), .A(PC_2_), .B(_3247__bF_buf2), .Q(_3251_) );
NA2X1 NA2X1_918 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2684_), .B(_3244__bF_buf3), .Q(_3252_) );
NA2X1 NA2X1_919 ( .gnd!(gnd!), .vdd!(vdd!), .A(PCU_ePC_2_), .B(CTRL_cu_pc_s4_bF_buf5), .Q(_3253_) );
AN31X1 AN31X1_92 ( .gnd!(gnd!), .vdd!(vdd!), .A(_3247__bF_buf2), .B(_3253_), .C(_3252_), .D(_3251_), .Q(_2641__2_) );
NO2X1 NO2X1_406 ( .gnd!(gnd!), .vdd!(vdd!), .A(PC_3_), .B(_3247__bF_buf1), .Q(_3254_) );
NA2X1 NA2X1_920 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2700_), .B(_3244__bF_buf2), .Q(_3255_) );
NA2X1 NA2X1_921 ( .gnd!(gnd!), .vdd!(vdd!), .A(PCU_ePC_3_), .B(CTRL_cu_pc_s4_bF_buf0), .Q(_3256_) );
AN31X1 AN31X1_93 ( .gnd!(gnd!), .vdd!(vdd!), .A(_3247__bF_buf1), .B(_3256_), .C(_3255_), .D(_3254_), .Q(_2641__3_) );
NA2X1 NA2X1_922 ( .gnd!(gnd!), .vdd!(vdd!), .A(_3246__bF_buf1), .B(PC_4_), .Q(_3257_) );
INX1 INX1_241 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_cu_pc_s0), .Q(_3258_) );
AND2X2 AND2X2_102 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_cu_pc_s0), .B(PCU_int_vec_4_), .Q(_3259_) );
AN211X1 AN211X1_24 ( .gnd!(gnd!), .vdd!(vdd!), .A(_3258_), .B(_2732_), .C(CTRL_cu_pc_s4_bF_buf2), .D(_3259_), .Q(_3260_) );
AND2X2 AND2X2_103 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2702_), .B(CTRL_cu_pc_s4_bF_buf2), .Q(_3261_) );
ON31X1 ON31X1_104 ( .gnd!(gnd!), .vdd!(vdd!), .A(_3246__bF_buf2), .B(_3261_), .C(_3260_), .D(_3257_), .Q(_2641__4_) );
NA2X1 NA2X1_923 ( .gnd!(gnd!), .vdd!(vdd!), .A(_3246__bF_buf1), .B(PC_5_), .Q(_3262_) );
AND2X2 AND2X2_104 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_cu_pc_s0), .B(PCU_int_vec_5_), .Q(_3263_) );
AN211X1 AN211X1_25 ( .gnd!(gnd!), .vdd!(vdd!), .A(_3258_), .B(_2744_), .C(CTRL_cu_pc_s4_bF_buf2), .D(_3263_), .Q(_3264_) );
AND2X2 AND2X2_105 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2734_), .B(CTRL_cu_pc_s4_bF_buf3), .Q(_3265_) );
ON31X1 ON31X1_105 ( .gnd!(gnd!), .vdd!(vdd!), .A(_3246__bF_buf1), .B(_3265_), .C(_3264_), .D(_3262_), .Q(_2641__5_) );
NA2X1 NA2X1_924 ( .gnd!(gnd!), .vdd!(vdd!), .A(_3246__bF_buf1), .B(PC_6_), .Q(_3266_) );
AND2X2 AND2X2_106 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_cu_pc_s0), .B(IRQ), .Q(_3267_) );
AN211X1 AN211X1_26 ( .gnd!(gnd!), .vdd!(vdd!), .A(_3258_), .B(_2760_), .C(CTRL_cu_pc_s4_bF_buf2), .D(_3267_), .Q(_3268_) );
AND2X2 AND2X2_107 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2746_), .B(CTRL_cu_pc_s4_bF_buf3), .Q(_3269_) );
ON31X1 ON31X1_106 ( .gnd!(gnd!), .vdd!(vdd!), .A(_3246__bF_buf1), .B(_3269_), .C(_3268_), .D(_3266_), .Q(_2641__6_) );
NO2X1 NO2X1_407 ( .gnd!(gnd!), .vdd!(vdd!), .A(PC_7_), .B(_3247__bF_buf0), .Q(_3270_) );
NA2X1 NA2X1_925 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2776_), .B(_3244__bF_buf3), .Q(_3271_) );
NA2X1 NA2X1_926 ( .gnd!(gnd!), .vdd!(vdd!), .A(PCU_ePC_7_), .B(CTRL_cu_pc_s4_bF_buf4), .Q(_3272_) );
AN31X1 AN31X1_94 ( .gnd!(gnd!), .vdd!(vdd!), .A(_3247__bF_buf4), .B(_3272_), .C(_3271_), .D(_3270_), .Q(_2641__7_) );
NO2X1 NO2X1_408 ( .gnd!(gnd!), .vdd!(vdd!), .A(PC_8_), .B(_3247__bF_buf1), .Q(_3273_) );
NA2X1 NA2X1_927 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2799_), .B(_3244__bF_buf2), .Q(_3274_) );
NA2X1 NA2X1_928 ( .gnd!(gnd!), .vdd!(vdd!), .A(PCU_ePC_8_), .B(CTRL_cu_pc_s4_bF_buf4), .Q(_3275_) );
AN31X1 AN31X1_95 ( .gnd!(gnd!), .vdd!(vdd!), .A(_3247__bF_buf1), .B(_3275_), .C(_3274_), .D(_3273_), .Q(_2641__8_) );
NO2X1 NO2X1_409 ( .gnd!(gnd!), .vdd!(vdd!), .A(PC_9_), .B(_3247__bF_buf4), .Q(_3276_) );
NA2X1 NA2X1_929 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2817_), .B(_3244__bF_buf1), .Q(_3277_) );
NA2X1 NA2X1_930 ( .gnd!(gnd!), .vdd!(vdd!), .A(PCU_ePC_9_), .B(CTRL_cu_pc_s4_bF_buf3), .Q(_3278_) );
AN31X1 AN31X1_96 ( .gnd!(gnd!), .vdd!(vdd!), .A(_3247__bF_buf4), .B(_3278_), .C(_3277_), .D(_3276_), .Q(_2641__9_) );
INX1 INX1_242 ( .gnd!(gnd!), .vdd!(vdd!), .A(_3244__bF_buf2), .Q(_3279_) );
NA3I1X1 NA3I1X1_130 ( .gnd!(gnd!), .vdd!(vdd!), .AN(_3279_), .B(_2834_), .C(_2833_), .Q(_3280_) );
AN21X1 AN21X1_193 ( .gnd!(gnd!), .vdd!(vdd!), .A(PCU_ePC_10_), .B(CTRL_cu_pc_s4_bF_buf4), .C(_3246__bF_buf3), .Q(_3281_) );
AN22X1 AN22X1_82 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2835_), .B(_3246__bF_buf4), .C(_3280_), .D(_3281_), .Q(_2641__10_) );
NO2X1 NO2X1_410 ( .gnd!(gnd!), .vdd!(vdd!), .A(PC_11_), .B(_3247__bF_buf2), .Q(_3282_) );
NA2X1 NA2X1_931 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2855_), .B(_3244__bF_buf4), .Q(_3283_) );
NA2X1 NA2X1_932 ( .gnd!(gnd!), .vdd!(vdd!), .A(PCU_ePC_11_), .B(CTRL_cu_pc_s4_bF_buf1), .Q(_3284_) );
AN31X1 AN31X1_97 ( .gnd!(gnd!), .vdd!(vdd!), .A(_3247__bF_buf3), .B(_3284_), .C(_3283_), .D(_3282_), .Q(_2641__11_) );
NO2X1 NO2X1_411 ( .gnd!(gnd!), .vdd!(vdd!), .A(PC_12_), .B(_3247__bF_buf3), .Q(_3285_) );
NA2X1 NA2X1_933 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2884_), .B(_3244__bF_buf4), .Q(_3286_) );
NA2X1 NA2X1_934 ( .gnd!(gnd!), .vdd!(vdd!), .A(PCU_ePC_12_), .B(CTRL_cu_pc_s4_bF_buf1), .Q(_3287_) );
AN31X1 AN31X1_98 ( .gnd!(gnd!), .vdd!(vdd!), .A(_3247__bF_buf3), .B(_3287_), .C(_3286_), .D(_3285_), .Q(_2641__12_) );
NO2X1 NO2X1_412 ( .gnd!(gnd!), .vdd!(vdd!), .A(PC_13_), .B(_3247__bF_buf3), .Q(_3288_) );
NA2X1 NA2X1_935 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2901_), .B(_3244__bF_buf4), .Q(_3289_) );
NA2X1 NA2X1_936 ( .gnd!(gnd!), .vdd!(vdd!), .A(PCU_ePC_13_), .B(CTRL_cu_pc_s4_bF_buf1), .Q(_3290_) );
AN31X1 AN31X1_99 ( .gnd!(gnd!), .vdd!(vdd!), .A(_3247__bF_buf3), .B(_3290_), .C(_3289_), .D(_3288_), .Q(_2641__13_) );
ON21X1 ON21X1_374 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2918_), .B(_2904_), .C(_3244__bF_buf1), .Q(_3291_) );
AN21X1 AN21X1_194 ( .gnd!(gnd!), .vdd!(vdd!), .A(PCU_ePC_14_), .B(CTRL_cu_pc_s4_bF_buf0), .C(_3246__bF_buf4), .Q(_3292_) );
AN22X1 AN22X1_83 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2910_), .B(_3246__bF_buf4), .C(_3291_), .D(_3292_), .Q(_2641__14_) );
NA2X1 NA2X1_937 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2933_), .B(_3244__bF_buf4), .Q(_3293_) );
AN21X1 AN21X1_195 ( .gnd!(gnd!), .vdd!(vdd!), .A(PCU_ePC_15_), .B(CTRL_cu_pc_s4_bF_buf1), .C(_3246__bF_buf2), .Q(_3294_) );
AN22X1 AN22X1_84 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2934_), .B(_3246__bF_buf2), .C(_3293_), .D(_3294_), .Q(_2641__15_) );
NA2X1 NA2X1_938 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2984_), .B(_3244__bF_buf0), .Q(_3295_) );
AN21X1 AN21X1_196 ( .gnd!(gnd!), .vdd!(vdd!), .A(PCU_ePC_16_), .B(CTRL_cu_pc_s4_bF_buf5), .C(_3246__bF_buf3), .Q(_3296_) );
AN22X1 AN22X1_85 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2962_), .B(_3246__bF_buf0), .C(_3295_), .D(_3296_), .Q(_2641__16_) );
NO2X1 NO2X1_413 ( .gnd!(gnd!), .vdd!(vdd!), .A(PC_17_), .B(_3247__bF_buf2), .Q(_3297_) );
NA2X1 NA2X1_939 ( .gnd!(gnd!), .vdd!(vdd!), .A(_2997_), .B(_3244__bF_buf3), .Q(_3298_) );
NA2X1 NA2X1_940 ( .gnd!(gnd!), .vdd!(vdd!), .A(PCU_ePC_17_), .B(CTRL_cu_pc_s4_bF_buf5), .Q(_3299_) );
AN31X1 AN31X1_100 ( .gnd!(gnd!), .vdd!(vdd!), .A(_3247__bF_buf2), .B(_3299_), .C(_3298_), .D(_3297_), .Q(_2641__17_) );
ON21X1 ON21X1_375 ( .gnd!(gnd!), .vdd!(vdd!), .A(_3013_), .B(_3000_), .C(_3244__bF_buf0), .Q(_3300_) );
AN21X1 AN21X1_197 ( .gnd!(gnd!), .vdd!(vdd!), .A(PCU_ePC_18_), .B(CTRL_cu_pc_s4_bF_buf4), .C(_3246__bF_buf3), .Q(_3301_) );
AN22X1 AN22X1_86 ( .gnd!(gnd!), .vdd!(vdd!), .A(_3008_), .B(_3246__bF_buf3), .C(_3300_), .D(_3301_), .Q(_2641__18_) );
NA2I1X1 NA2I1X1_142 ( .gnd!(gnd!), .vdd!(vdd!), .AN(_3030_), .B(_3244__bF_buf0), .Q(_3302_) );
AN21X1 AN21X1_198 ( .gnd!(gnd!), .vdd!(vdd!), .A(PCU_ePC_19_), .B(CTRL_cu_pc_s4_bF_buf5), .C(_3246__bF_buf0), .Q(_3303_) );
AN22X1 AN22X1_87 ( .gnd!(gnd!), .vdd!(vdd!), .A(_3016_), .B(_3246__bF_buf0), .C(_3302_), .D(_3303_), .Q(_2641__19_) );
NA2X1 NA2X1_941 ( .gnd!(gnd!), .vdd!(vdd!), .A(_3048_), .B(_3244__bF_buf0), .Q(_3304_) );
AN21X1 AN21X1_199 ( .gnd!(gnd!), .vdd!(vdd!), .A(PCU_ePC_20_), .B(CTRL_cu_pc_s4_bF_buf5), .C(_3246__bF_buf3), .Q(_3305_) );
AN22X1 AN22X1_88 ( .gnd!(gnd!), .vdd!(vdd!), .A(_3040_), .B(_3246__bF_buf0), .C(_3304_), .D(_3305_), .Q(_2641__20_) );
NA2X1 NA2X1_942 ( .gnd!(gnd!), .vdd!(vdd!), .A(_3075_), .B(_3244__bF_buf0), .Q(_3306_) );
AN21X1 AN21X1_200 ( .gnd!(gnd!), .vdd!(vdd!), .A(PCU_ePC_21_), .B(CTRL_cu_pc_s4_bF_buf5), .C(_3246__bF_buf0), .Q(_3307_) );
AN22X1 AN22X1_89 ( .gnd!(gnd!), .vdd!(vdd!), .A(_3062_), .B(_3246__bF_buf0), .C(_3306_), .D(_3307_), .Q(_2641__21_) );
NO2X1 NO2X1_414 ( .gnd!(gnd!), .vdd!(vdd!), .A(PC_22_), .B(_3247__bF_buf2), .Q(_3308_) );
ON21X1 ON21X1_376 ( .gnd!(gnd!), .vdd!(vdd!), .A(_3091_), .B(_3078_), .C(_3244__bF_buf3), .Q(_3309_) );
NA2X1 NA2X1_943 ( .gnd!(gnd!), .vdd!(vdd!), .A(PCU_ePC_22_), .B(CTRL_cu_pc_s4_bF_buf5), .Q(_3310_) );
AN31X1 AN31X1_101 ( .gnd!(gnd!), .vdd!(vdd!), .A(_3247__bF_buf0), .B(_3310_), .C(_3309_), .D(_3308_), .Q(_2641__22_) );
NA3I1X1 NA3I1X1_131 ( .gnd!(gnd!), .vdd!(vdd!), .AN(_3279_), .B(_3095_), .C(_3107_), .Q(_3311_) );
AN21X1 AN21X1_201 ( .gnd!(gnd!), .vdd!(vdd!), .A(PCU_ePC_23_), .B(CTRL_cu_pc_s4_bF_buf4), .C(_3246__bF_buf3), .Q(_3312_) );
AN22X1 AN22X1_90 ( .gnd!(gnd!), .vdd!(vdd!), .A(_3097_), .B(_3246__bF_buf3), .C(_3311_), .D(_3312_), .Q(_2641__23_) );
NO2X1 NO2X1_415 ( .gnd!(gnd!), .vdd!(vdd!), .A(PC_24_), .B(_3247__bF_buf0), .Q(_3313_) );
NA2X1 NA2X1_944 ( .gnd!(gnd!), .vdd!(vdd!), .A(_3135_), .B(_3244__bF_buf3), .Q(_3314_) );
NA2X1 NA2X1_945 ( .gnd!(gnd!), .vdd!(vdd!), .A(PCU_ePC_24_), .B(CTRL_cu_pc_s4_bF_buf3), .Q(_3315_) );
AN31X1 AN31X1_102 ( .gnd!(gnd!), .vdd!(vdd!), .A(_3247__bF_buf0), .B(_3315_), .C(_3314_), .D(_3313_), .Q(_2641__24_) );
NO2X1 NO2X1_416 ( .gnd!(gnd!), .vdd!(vdd!), .A(PC_25_), .B(_3247__bF_buf1), .Q(_3316_) );
NA2X1 NA2X1_946 ( .gnd!(gnd!), .vdd!(vdd!), .A(_3149_), .B(_3244__bF_buf2), .Q(_3317_) );
NA2X1 NA2X1_947 ( .gnd!(gnd!), .vdd!(vdd!), .A(PCU_ePC_25_), .B(CTRL_cu_pc_s4_bF_buf0), .Q(_3318_) );
AN31X1 AN31X1_103 ( .gnd!(gnd!), .vdd!(vdd!), .A(_3247__bF_buf1), .B(_3318_), .C(_3317_), .D(_3316_), .Q(_2641__25_) );
NO2X1 NO2X1_417 ( .gnd!(gnd!), .vdd!(vdd!), .A(PC_26_), .B(_3247__bF_buf0), .Q(_3319_) );
ON21X1 ON21X1_377 ( .gnd!(gnd!), .vdd!(vdd!), .A(_3162_), .B(_3152_), .C(_3244__bF_buf3), .Q(_3320_) );
NA2X1 NA2X1_948 ( .gnd!(gnd!), .vdd!(vdd!), .A(PCU_ePC_26_), .B(CTRL_cu_pc_s4_bF_buf4), .Q(_3321_) );
AN31X1 AN31X1_104 ( .gnd!(gnd!), .vdd!(vdd!), .A(_3247__bF_buf0), .B(_3321_), .C(_3320_), .D(_3319_), .Q(_2641__26_) );
NA3I1X1 NA3I1X1_132 ( .gnd!(gnd!), .vdd!(vdd!), .AN(_3279_), .B(_3166_), .C(_3174_), .Q(_3322_) );
AN21X1 AN21X1_202 ( .gnd!(gnd!), .vdd!(vdd!), .A(PCU_ePC_27_), .B(CTRL_cu_pc_s4_bF_buf0), .C(_3246__bF_buf4), .Q(_3323_) );
AN22X1 AN22X1_91 ( .gnd!(gnd!), .vdd!(vdd!), .A(_3175_), .B(_3246__bF_buf4), .C(_3322_), .D(_3323_), .Q(_2641__27_) );
NO2X1 NO2X1_418 ( .gnd!(gnd!), .vdd!(vdd!), .A(PC_28_), .B(_3247__bF_buf4), .Q(_3324_) );
NA2X1 NA2X1_949 ( .gnd!(gnd!), .vdd!(vdd!), .A(_3196_), .B(_3244__bF_buf2), .Q(_3325_) );
NA2X1 NA2X1_950 ( .gnd!(gnd!), .vdd!(vdd!), .A(PCU_ePC_28_), .B(CTRL_cu_pc_s4_bF_buf0), .Q(_3326_) );
AN31X1 AN31X1_105 ( .gnd!(gnd!), .vdd!(vdd!), .A(_3247__bF_buf4), .B(_3326_), .C(_3325_), .D(_3324_), .Q(_2641__28_) );
NA2X1 NA2X1_951 ( .gnd!(gnd!), .vdd!(vdd!), .A(_3210_), .B(_3244__bF_buf4), .Q(_3327_) );
AN21X1 AN21X1_203 ( .gnd!(gnd!), .vdd!(vdd!), .A(PCU_ePC_29_), .B(CTRL_cu_pc_s4_bF_buf1), .C(_3246__bF_buf2), .Q(_3328_) );
AN22X1 AN22X1_92 ( .gnd!(gnd!), .vdd!(vdd!), .A(_3211_), .B(_3246__bF_buf2), .C(_3327_), .D(_3328_), .Q(_2641__29_) );
NO2X1 NO2X1_419 ( .gnd!(gnd!), .vdd!(vdd!), .A(PC_30_), .B(_3247__bF_buf4), .Q(_3329_) );
ON21X1 ON21X1_378 ( .gnd!(gnd!), .vdd!(vdd!), .A(_3228_), .B(CTRL_IDEC1_cu_jalr_inst_bF_buf0), .C(_3229_), .Q(_3330_) );
NA2X1 NA2X1_952 ( .gnd!(gnd!), .vdd!(vdd!), .A(_3330_), .B(_3244__bF_buf1), .Q(_3331_) );
NA2X1 NA2X1_953 ( .gnd!(gnd!), .vdd!(vdd!), .A(PCU_ePC_30_), .B(CTRL_cu_pc_s4_bF_buf0), .Q(_3332_) );
AN31X1 AN31X1_106 ( .gnd!(gnd!), .vdd!(vdd!), .A(_3247__bF_buf4), .B(_3332_), .C(_3331_), .D(_3329_), .Q(_2641__30_) );
INX1 INX1_243 ( .gnd!(gnd!), .vdd!(vdd!), .A(PC_31_), .Q(_3333_) );
OA211X4 OA211X4_3 ( .gnd!(gnd!), .vdd!(vdd!), .A(_3216_), .B(_3220_), .C(_3221_), .D(_3237_), .Q(_3334_) );
AN21X1 AN21X1_204 ( .gnd!(gnd!), .vdd!(vdd!), .A(_3227_), .B(_3221_), .C(_3237_), .Q(_3335_) );
NA2X1 NA2X1_954 ( .gnd!(gnd!), .vdd!(vdd!), .A(_3240_), .B(CTRL_IDEC1_cu_jalr_inst_bF_buf3), .Q(_3336_) );
ON311X1 ON311X1_18 ( .gnd!(gnd!), .vdd!(vdd!), .A(CTRL_IDEC1_cu_jalr_inst_bF_buf3), .B(_3334_), .C(_3335_), .D(_3336_), .E(_3244__bF_buf1), .Q(_3337_) );
AN21X1 AN21X1_205 ( .gnd!(gnd!), .vdd!(vdd!), .A(PCU_ePC_31_), .B(CTRL_cu_pc_s4_bF_buf3), .C(_3246__bF_buf4), .Q(_3338_) );
AN22X1 AN22X1_93 ( .gnd!(gnd!), .vdd!(vdd!), .A(_3333_), .B(_3246__bF_buf4), .C(_3337_), .D(_3338_), .Q(_2641__31_) );
INX3 INX3_9 ( .gnd!(gnd!), .vdd!(vdd!), .A(rst), .Q(_3117_) );
DFRRQX1 DFRRQX1_184 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf0), .D(_2642__0_), .Q(PCU_ePC_0_), .RN(_3117__bF_buf3) );
DFRRQX1 DFRRQX1_185 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf18), .D(_2642__1_), .Q(PCU_ePC_1_), .RN(_3117__bF_buf4) );
DFRRQX1 DFRRQX1_186 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf35), .D(_2642__2_), .Q(PCU_ePC_2_), .RN(_3117__bF_buf0) );
DFRRQX1 DFRRQX1_187 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf38), .D(_2642__3_), .Q(PCU_ePC_3_), .RN(_3117__bF_buf5) );
DFRRQX1 DFRRQX1_188 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf18), .D(_2642__4_), .Q(PCU_ePC_4_), .RN(_3117__bF_buf4) );
DFRRQX1 DFRRQX1_189 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf0), .D(_2642__5_), .Q(PCU_ePC_5_), .RN(_3117__bF_buf3) );
DFRRQX1 DFRRQX1_190 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf0), .D(_2642__6_), .Q(PCU_ePC_6_), .RN(_3117__bF_buf3) );
DFRRQX1 DFRRQX1_191 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf3), .D(_2642__7_), .Q(PCU_ePC_7_), .RN(_3117__bF_buf2) );
DFRRQX1 DFRRQX1_192 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf15), .D(_2642__8_), .Q(PCU_ePC_8_), .RN(_3117__bF_buf2) );
DFRRQX1 DFRRQX1_193 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf51), .D(_2642__9_), .Q(PCU_ePC_9_), .RN(_3117__bF_buf1) );
DFRRQX1 DFRRQX1_194 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf38), .D(_2642__10_), .Q(PCU_ePC_10_), .RN(_3117__bF_buf5) );
DFRRQX1 DFRRQX1_195 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf35), .D(_2642__11_), .Q(PCU_ePC_11_), .RN(_3117__bF_buf0) );
DFRRQX1 DFRRQX1_196 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf35), .D(_2642__12_), .Q(PCU_ePC_12_), .RN(_3117__bF_buf4) );
DFRRQX1 DFRRQX1_197 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf18), .D(_2642__13_), .Q(PCU_ePC_13_), .RN(_3117__bF_buf4) );
DFRRQX1 DFRRQX1_198 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf51), .D(_2642__14_), .Q(PCU_ePC_14_), .RN(_3117__bF_buf1) );
DFRRQX1 DFRRQX1_199 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf52), .D(_2642__15_), .Q(PCU_ePC_15_), .RN(_3117__bF_buf4) );
DFRRQX1 DFRRQX1_200 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf25), .D(_2642__16_), .Q(PCU_ePC_16_), .RN(_3117__bF_buf6) );
DFRRQX1 DFRRQX1_201 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf3), .D(_2642__17_), .Q(PCU_ePC_17_), .RN(_3117__bF_buf2) );
DFRRQX1 DFRRQX1_202 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf15), .D(_2642__18_), .Q(PCU_ePC_18_), .RN(_3117__bF_buf5) );
DFRRQX1 DFRRQX1_203 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf25), .D(_2642__19_), .Q(PCU_ePC_19_), .RN(_3117__bF_buf6) );
DFRRQX1 DFRRQX1_204 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf3), .D(_2642__20_), .Q(PCU_ePC_20_), .RN(_3117__bF_buf2) );
DFRRQX1 DFRRQX1_205 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf25), .D(_2642__21_), .Q(PCU_ePC_21_), .RN(_3117__bF_buf6) );
DFRRQX1 DFRRQX1_206 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf3), .D(_2642__22_), .Q(PCU_ePC_22_), .RN(_3117__bF_buf2) );
DFRRQX1 DFRRQX1_207 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf25), .D(_2642__23_), .Q(PCU_ePC_23_), .RN(_3117__bF_buf6) );
DFRRQX1 DFRRQX1_208 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf49), .D(_2642__24_), .Q(PCU_ePC_24_), .RN(_3117__bF_buf3) );
DFRRQX1 DFRRQX1_209 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf15), .D(_2642__25_), .Q(PCU_ePC_25_), .RN(_3117__bF_buf7) );
DFRRQX1 DFRRQX1_210 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf49), .D(_2642__26_), .Q(PCU_ePC_26_), .RN(_3117__bF_buf2) );
DFRRQX1 DFRRQX1_211 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf49), .D(_2642__27_), .Q(PCU_ePC_27_), .RN(_3117__bF_buf7) );
DFRRQX1 DFRRQX1_212 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf49), .D(_2642__28_), .Q(PCU_ePC_28_), .RN(_3117__bF_buf7) );
DFRRQX1 DFRRQX1_213 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf18), .D(_2642__29_), .Q(PCU_ePC_29_), .RN(_3117__bF_buf4) );
DFRRQX1 DFRRQX1_214 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf38), .D(_2642__30_), .Q(PCU_ePC_30_), .RN(_3117__bF_buf1) );
DFRRQX1 DFRRQX1_215 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf51), .D(_2642__31_), .Q(PCU_ePC_31_), .RN(_3117__bF_buf1) );
DFRRQX1 DFRRQX1_216 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf51), .D(_2641__0_), .Q(PC_0_), .RN(_3117__bF_buf3) );
DFRRQX1 DFRRQX1_217 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf35), .D(_2641__1_), .Q(PC_1_), .RN(_3117__bF_buf4) );
DFRRQX1 DFRRQX1_218 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf35), .D(_2641__2_), .Q(PC_2_), .RN(_3117__bF_buf0) );
DFRRQX1 DFRRQX1_219 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf38), .D(_2641__3_), .Q(PC_3_), .RN(_3117__bF_buf7) );
DFRRQX1 DFRRQX1_220 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf0), .D(_2641__4_), .Q(PC_4_), .RN(_3117__bF_buf0) );
DFRRQX1 DFRRQX1_221 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf51), .D(_2641__5_), .Q(PC_5_), .RN(_3117__bF_buf3) );
DFRRQX1 DFRRQX1_222 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf0), .D(_2641__6_), .Q(PC_6_), .RN(_3117__bF_buf3) );
DFRRQX1 DFRRQX1_223 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf3), .D(_2641__7_), .Q(PC_7_), .RN(_3117__bF_buf2) );
DFRRQX1 DFRRQX1_224 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf15), .D(_2641__8_), .Q(PC_8_), .RN(_3117__bF_buf5) );
DFRRQX1 DFRRQX1_225 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf49), .D(_2641__9_), .Q(PC_9_), .RN(_3117__bF_buf1) );
DFRRQX1 DFRRQX1_226 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf38), .D(_2641__10_), .Q(PC_10_), .RN(_3117__bF_buf5) );
DFRRQX1 DFRRQX1_227 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf35), .D(_2641__11_), .Q(PC_11_), .RN(_3117__bF_buf0) );
DFRRQX1 DFRRQX1_228 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf18), .D(_2641__12_), .Q(PC_12_), .RN(_3117__bF_buf4) );
DFRRQX1 DFRRQX1_229 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf35), .D(_2641__13_), .Q(PC_13_), .RN(_3117__bF_buf0) );
DFRRQX1 DFRRQX1_230 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf38), .D(_2641__14_), .Q(PC_14_), .RN(_3117__bF_buf1) );
DFRRQX1 DFRRQX1_231 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf49), .D(_2641__15_), .Q(PC_15_), .RN(_3117__bF_buf3) );
DFRRQX1 DFRRQX1_232 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf25), .D(_2641__16_), .Q(PC_16_), .RN(_3117__bF_buf6) );
DFRRQX1 DFRRQX1_233 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf3), .D(_2641__17_), .Q(PC_17_), .RN(_3117__bF_buf2) );
DFRRQX1 DFRRQX1_234 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf15), .D(_2641__18_), .Q(PC_18_), .RN(_3117__bF_buf5) );
DFRRQX1 DFRRQX1_235 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf3), .D(_2641__19_), .Q(PC_19_), .RN(_3117__bF_buf6) );
DFRRQX1 DFRRQX1_236 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf25), .D(_2641__20_), .Q(PC_20_), .RN(_3117__bF_buf6) );
DFRRQX1 DFRRQX1_237 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf25), .D(_2641__21_), .Q(PC_21_), .RN(_3117__bF_buf6) );
DFRRQX1 DFRRQX1_238 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf35), .D(_2641__22_), .Q(PC_22_), .RN(_3117__bF_buf0) );
DFRRQX1 DFRRQX1_239 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf15), .D(_2641__23_), .Q(PC_23_), .RN(_3117__bF_buf5) );
DFRRQX1 DFRRQX1_240 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf49), .D(_2641__24_), .Q(PC_24_), .RN(_3117__bF_buf7) );
DFRRQX1 DFRRQX1_241 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf15), .D(_2641__25_), .Q(PC_25_), .RN(_3117__bF_buf7) );
DFRRQX1 DFRRQX1_242 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf49), .D(_2641__26_), .Q(PC_26_), .RN(_3117__bF_buf7) );
DFRRQX1 DFRRQX1_243 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf38), .D(_2641__27_), .Q(PC_27_), .RN(_3117__bF_buf5) );
DFRRQX1 DFRRQX1_244 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf38), .D(_2641__28_), .Q(PC_28_), .RN(_3117__bF_buf7) );
DFRRQX1 DFRRQX1_245 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf52), .D(_2641__29_), .Q(PC_29_), .RN(_3117__bF_buf0) );
DFRRQX1 DFRRQX1_246 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf51), .D(_2641__30_), .Q(PC_30_), .RN(_3117__bF_buf1) );
DFRRQX1 DFRRQX1_247 ( .gnd!(gnd!), .vdd!(vdd!), .C(clk_bF_buf51), .D(_2641__31_), .Q(PC_31_), .RN(_3117__bF_buf1) );
endmodule
