// file: memory.v
// author: @shalan


//`define _MEMDISP_ 	0

//MM IO
`define    MMAP_PRINT	32'h80000000
`define    LOGCAPH	12 

module rv32i_mem_ctrl (baddr, addr_targ, bsz, bdi, mdi, mcs, bdo, mdo);
    input[1:0] baddr;
    input addr_targ;
    input[1:0] bsz;
    input[31:0] bdi, mdo;
    
    output [31:0] bdo;
    output reg [31:0] mdi;
    output reg [3:0] mcs;
    
    reg [31:0] bdo_reg;
    
    wire szB=(bsz==2'b0);
    wire szH=(bsz==2'b01);
    wire szW=(bsz==2'b10);

    always @ * begin
    (* full_case *)
        (* parallel_case *)
        case ({baddr, szB, szH, szW})
            5'b00_001: begin mdi = bdi; mcs=4'b1111; end

            5'b00_010: begin mdi = bdi; mcs=4'b0011; end
            5'b10_010: begin mdi = bdi << 16; mcs=4'b1100; end

            5'b00_100: begin mdi = bdi; mcs=4'b0001; end
            5'b01_100: begin mdi = bdi << 8; mcs=4'b0010; end
            5'b10_100: begin mdi = bdi << 16; mcs=4'b0100; end
            5'b11_100: begin mdi = bdi << 24; mcs=4'b1000; end
        endcase

    end

    always @ * begin
    (* full_case *)
        (* parallel_case *)
        case ({baddr, szB, szH, szW})
            5'b00_001: bdo_reg = mdo;

            5'b00_010: bdo_reg = mdo;
            5'b10_010: bdo_reg = mdo >> 16;

            5'b00_100: bdo_reg = mdo;
            5'b01_100: bdo_reg = mdo >> 8;
            5'b10_100: bdo_reg = mdo >> 16;
            5'b11_100: bdo_reg = mdo >> 24;
        endcase
    end
    
    assign bdo = addr_targ? bdo_reg : 32'hZZZZZZZZ;

endmodule


module memory #(parameter capH = 1024) (input clk, input[31:0] bdi, baddr, output[31:0] bdo, input bwr, input[1:0] bsz );
    reg[7:0] bank0[capH-1:0];
    reg[7:0] bank1[capH-1:0];
    reg[7:0] bank2[capH-1:0];
    reg[7:0] bank3[capH-1:0];

    wire[31:0] mdo, mdi;
    wire[3:0] mcs;
    wire mwr;
    wire addr_targ =  (baddr[31:16] == 16'b0); //optimize using LOGCAPH 
    
    rv32i_mem_ctrl MCTRL (.baddr(baddr[1:0]), .addr_targ(addr_targ), .bsz(bsz), .bdi(bdi), .mdi(mdi), .mcs(mcs), .bdo(bdo), .mdo(mdo));

    assign mdo = {bank3[baddr[`LOGCAPH-1:2]],bank2[baddr[`LOGCAPH-1:2]],bank1[baddr[`LOGCAPH-1:2]],bank0[baddr[`LOGCAPH-1:2]]};
    assign mwr = bwr & addr_targ; 
    always @(posedge clk) begin
	    if (mwr) begin
				if(mcs[0]) bank0[baddr[`LOGCAPH-1:2]] <= mdi[7:0];
				if(mcs[1]) bank1[baddr[`LOGCAPH-1:2]] <= mdi[15:8];
				if(mcs[2]) bank2[baddr[`LOGCAPH-1:2]] <= mdi[23:16];
				if(mcs[3]) bank3[baddr[`LOGCAPH-1:2]] <= mdi[31:24];
	    end
    end


    //fpga only; rewrite using readmemh for each bank (change b2h_fpga.py to produce 4 files)
    initial begin   
    {bank3[0], bank2[0], bank1[0], bank0[0]} = 32'h00401073;
    {bank3[1], bank2[1], bank1[1], bank0[1]} = 32'h00000213;
    {bank3[2], bank2[2], bank1[2], bank0[2]} = 32'hc0121073;
    {bank3[3], bank2[3], bank1[3], bank0[3]} = 32'h0740006f;
    {bank3[4], bank2[4], bank1[4], bank0[4]} = 32'h00000013;
    {bank3[5], bank2[5], bank1[5], bank0[5]} = 32'h00200073;
    {bank3[6], bank2[6], bank1[6], bank0[6]} = 32'h00000000;
    {bank3[7], bank2[7], bank1[7], bank0[7]} = 32'h00000000;
    {bank3[8], bank2[8], bank1[8], bank0[8]} = 32'h00000013;
    {bank3[9], bank2[9], bank1[9], bank0[9]} = 32'h00200073;
    {bank3[10], bank2[10], bank1[10], bank0[10]} = 32'h00000000;
    {bank3[11], bank2[11], bank1[11], bank0[11]} = 32'h00000000;
    {bank3[12], bank2[12], bank1[12], bank0[12]} = 32'h01e00213;
    {bank3[13], bank2[13], bank1[13], bank0[13]} = 32'hc0121073;
    {bank3[14], bank2[14], bank1[14], bank0[14]} = 32'h00200073;
    {bank3[15], bank2[15], bank1[15], bank0[15]} = 32'h00000000;
    {bank3[16], bank2[16], bank1[16], bank0[16]} = 32'h0700006f;
    {bank3[17], bank2[17], bank1[17], bank0[17]} = 32'h0700006f;
    {bank3[18], bank2[18], bank1[18], bank0[18]} = 32'h0700006f;
    {bank3[19], bank2[19], bank1[19], bank0[19]} = 32'h0700006f;
    {bank3[20], bank2[20], bank1[20], bank0[20]} = 32'h0700006f;
    {bank3[21], bank2[21], bank1[21], bank0[21]} = 32'h0700006f;
    {bank3[22], bank2[22], bank1[22], bank0[22]} = 32'h0700006f;
    {bank3[23], bank2[23], bank1[23], bank0[23]} = 32'h0700006f;
    {bank3[24], bank2[24], bank1[24], bank0[24]} = 32'h0700006f;
    {bank3[25], bank2[25], bank1[25], bank0[25]} = 32'h0700006f;
    {bank3[26], bank2[26], bank1[26], bank0[26]} = 32'h0700006f;
    {bank3[27], bank2[27], bank1[27], bank0[27]} = 32'h0700006f;
    {bank3[28], bank2[28], bank1[28], bank0[28]} = 32'h0700006f;
    {bank3[29], bank2[29], bank1[29], bank0[29]} = 32'h0700006f;
    {bank3[30], bank2[30], bank1[30], bank0[30]} = 32'h0700006f;
    {bank3[31], bank2[31], bank1[31], bank0[31]} = 32'h0700006f;
    {bank3[32], bank2[32], bank1[32], bank0[32]} = 32'h00700213;
    {bank3[33], bank2[33], bank1[33], bank0[33]} = 32'h00421073;
    {bank3[34], bank2[34], bank1[34], bank0[34]} = 32'h00000137;
    {bank3[35], bank2[35], bank1[35], bank0[35]} = 32'h00010113;
    {bank3[36], bank2[36], bank1[36], bank0[36]} = 32'h00c000ef;
    {bank3[37], bank2[37], bank1[37], bank0[37]} = 32'h00a00893;
    {bank3[38], bank2[38], bank1[38], bank0[38]} = 32'h00000073;
    {bank3[39], bank2[39], bank1[39], bank0[39]} = 32'h800002b7;
    {bank3[40], bank2[40], bank1[40], bank0[40]} = 32'h0012a403;
    {bank3[41], bank2[41], bank1[41], bank0[41]} = 32'h00147313;
    {bank3[42], bank2[42], bank1[42], bank0[42]} = 32'hfe030ce3;
    {bank3[43], bank2[43], bank1[43], bank0[43]} = 32'h00008067;
    {bank3[44], bank2[44], bank1[44], bank0[44]} = 32'h00200073;
    {bank3[45], bank2[45], bank1[45], bank0[45]} = 32'h00200073;
    {bank3[46], bank2[46], bank1[46], bank0[46]} = 32'h00200073;
    {bank3[47], bank2[47], bank1[47], bank0[47]} = 32'h00200073;
    {bank3[48], bank2[48], bank1[48], bank0[48]} = 32'h00200073;
    {bank3[49], bank2[49], bank1[49], bank0[49]} = 32'h00200073;
    {bank3[50], bank2[50], bank1[50], bank0[50]} = 32'h00200073;
    {bank3[51], bank2[51], bank1[51], bank0[51]} = 32'h00200073;
    {bank3[52], bank2[52], bank1[52], bank0[52]} = 32'h00200073;
    {bank3[53], bank2[53], bank1[53], bank0[53]} = 32'h00200073;
    {bank3[54], bank2[54], bank1[54], bank0[54]} = 32'h00200073;
    {bank3[55], bank2[55], bank1[55], bank0[55]} = 32'h00200073;
    {bank3[56], bank2[56], bank1[56], bank0[56]} = 32'h00200073;
    {bank3[57], bank2[57], bank1[57], bank0[57]} = 32'h00200073;
    {bank3[58], bank2[58], bank1[58], bank0[58]} = 32'h00200073;
    {bank3[59], bank2[59], bank1[59], bank0[59]} = 32'h00200073;
    {bank3[60], bank2[60], bank1[60], bank0[60]} = 32'h0;
    {bank3[61], bank2[61], bank1[61], bank0[61]} = 32'h0;
    {bank3[62], bank2[62], bank1[62], bank0[62]} = 32'h0;
    {bank3[63], bank2[63], bank1[63], bank0[63]} = 32'h0;
    {bank3[64], bank2[64], bank1[64], bank0[64]} = 32'h0;
    {bank3[65], bank2[65], bank1[65], bank0[65]} = 32'h0;
    {bank3[66], bank2[66], bank1[66], bank0[66]} = 32'h0;
    {bank3[67], bank2[67], bank1[67], bank0[67]} = 32'h0;
    {bank3[68], bank2[68], bank1[68], bank0[68]} = 32'h0;
    {bank3[69], bank2[69], bank1[69], bank0[69]} = 32'h0;
    {bank3[70], bank2[70], bank1[70], bank0[70]} = 32'h0;
    {bank3[71], bank2[71], bank1[71], bank0[71]} = 32'h0;
    {bank3[72], bank2[72], bank1[72], bank0[72]} = 32'h0;
    {bank3[73], bank2[73], bank1[73], bank0[73]} = 32'h0;
    {bank3[74], bank2[74], bank1[74], bank0[74]} = 32'h0;
    {bank3[75], bank2[75], bank1[75], bank0[75]} = 32'h0;
    {bank3[76], bank2[76], bank1[76], bank0[76]} = 32'h0;
    {bank3[77], bank2[77], bank1[77], bank0[77]} = 32'h0;
    {bank3[78], bank2[78], bank1[78], bank0[78]} = 32'h0;
    {bank3[79], bank2[79], bank1[79], bank0[79]} = 32'h0;
    {bank3[80], bank2[80], bank1[80], bank0[80]} = 32'h0;
    {bank3[81], bank2[81], bank1[81], bank0[81]} = 32'h0;
    {bank3[82], bank2[82], bank1[82], bank0[82]} = 32'h0;
    {bank3[83], bank2[83], bank1[83], bank0[83]} = 32'h0;
    {bank3[84], bank2[84], bank1[84], bank0[84]} = 32'h0;
    {bank3[85], bank2[85], bank1[85], bank0[85]} = 32'h0;
    {bank3[86], bank2[86], bank1[86], bank0[86]} = 32'h0;
    {bank3[87], bank2[87], bank1[87], bank0[87]} = 32'h0;
    {bank3[88], bank2[88], bank1[88], bank0[88]} = 32'h0;
    {bank3[89], bank2[89], bank1[89], bank0[89]} = 32'h0;
    {bank3[90], bank2[90], bank1[90], bank0[90]} = 32'h0;
    {bank3[91], bank2[91], bank1[91], bank0[91]} = 32'h0;
    {bank3[92], bank2[92], bank1[92], bank0[92]} = 32'h0;
    {bank3[93], bank2[93], bank1[93], bank0[93]} = 32'h0;
    {bank3[94], bank2[94], bank1[94], bank0[94]} = 32'h0;
    {bank3[95], bank2[95], bank1[95], bank0[95]} = 32'h0;
    {bank3[96], bank2[96], bank1[96], bank0[96]} = 32'h0;
    {bank3[97], bank2[97], bank1[97], bank0[97]} = 32'h0;
    {bank3[98], bank2[98], bank1[98], bank0[98]} = 32'h0;
    {bank3[99], bank2[99], bank1[99], bank0[99]} = 32'h0;
    {bank3[100], bank2[100], bank1[100], bank0[100]} = 32'h0;
    {bank3[101], bank2[101], bank1[101], bank0[101]} = 32'h0;
    {bank3[102], bank2[102], bank1[102], bank0[102]} = 32'h0;
    {bank3[103], bank2[103], bank1[103], bank0[103]} = 32'h0;
    {bank3[104], bank2[104], bank1[104], bank0[104]} = 32'h0;
    {bank3[105], bank2[105], bank1[105], bank0[105]} = 32'h0;
    {bank3[106], bank2[106], bank1[106], bank0[106]} = 32'h0;
    {bank3[107], bank2[107], bank1[107], bank0[107]} = 32'h0;
    {bank3[108], bank2[108], bank1[108], bank0[108]} = 32'h0;
    {bank3[109], bank2[109], bank1[109], bank0[109]} = 32'h0;
    {bank3[110], bank2[110], bank1[110], bank0[110]} = 32'h0;
    {bank3[111], bank2[111], bank1[111], bank0[111]} = 32'h0;
    {bank3[112], bank2[112], bank1[112], bank0[112]} = 32'h0;
    {bank3[113], bank2[113], bank1[113], bank0[113]} = 32'h0;
    {bank3[114], bank2[114], bank1[114], bank0[114]} = 32'h0;
    {bank3[115], bank2[115], bank1[115], bank0[115]} = 32'h0;
    {bank3[116], bank2[116], bank1[116], bank0[116]} = 32'h0;
    {bank3[117], bank2[117], bank1[117], bank0[117]} = 32'h0;
    {bank3[118], bank2[118], bank1[118], bank0[118]} = 32'h0;
    {bank3[119], bank2[119], bank1[119], bank0[119]} = 32'h0;
    {bank3[120], bank2[120], bank1[120], bank0[120]} = 32'h0;
    {bank3[121], bank2[121], bank1[121], bank0[121]} = 32'h0;
    {bank3[122], bank2[122], bank1[122], bank0[122]} = 32'h0;
    {bank3[123], bank2[123], bank1[123], bank0[123]} = 32'h0;
    {bank3[124], bank2[124], bank1[124], bank0[124]} = 32'h0;
    {bank3[125], bank2[125], bank1[125], bank0[125]} = 32'h0;
    {bank3[126], bank2[126], bank1[126], bank0[126]} = 32'h0;
    {bank3[127], bank2[127], bank1[127], bank0[127]} = 32'h0;
    {bank3[128], bank2[128], bank1[128], bank0[128]} = 32'h0;
    {bank3[129], bank2[129], bank1[129], bank0[129]} = 32'h0;
    {bank3[130], bank2[130], bank1[130], bank0[130]} = 32'h0;
    {bank3[131], bank2[131], bank1[131], bank0[131]} = 32'h0;
    {bank3[132], bank2[132], bank1[132], bank0[132]} = 32'h0;
    {bank3[133], bank2[133], bank1[133], bank0[133]} = 32'h0;
    {bank3[134], bank2[134], bank1[134], bank0[134]} = 32'h0;
    {bank3[135], bank2[135], bank1[135], bank0[135]} = 32'h0;
    {bank3[136], bank2[136], bank1[136], bank0[136]} = 32'h0;
    {bank3[137], bank2[137], bank1[137], bank0[137]} = 32'h0;
    {bank3[138], bank2[138], bank1[138], bank0[138]} = 32'h0;
    {bank3[139], bank2[139], bank1[139], bank0[139]} = 32'h0;
    {bank3[140], bank2[140], bank1[140], bank0[140]} = 32'h0;
    {bank3[141], bank2[141], bank1[141], bank0[141]} = 32'h0;
    {bank3[142], bank2[142], bank1[142], bank0[142]} = 32'h0;
    {bank3[143], bank2[143], bank1[143], bank0[143]} = 32'h0;
    {bank3[144], bank2[144], bank1[144], bank0[144]} = 32'h0;
    {bank3[145], bank2[145], bank1[145], bank0[145]} = 32'h0;
    {bank3[146], bank2[146], bank1[146], bank0[146]} = 32'h0;
    {bank3[147], bank2[147], bank1[147], bank0[147]} = 32'h0;
    {bank3[148], bank2[148], bank1[148], bank0[148]} = 32'h0;
    {bank3[149], bank2[149], bank1[149], bank0[149]} = 32'h0;
    {bank3[150], bank2[150], bank1[150], bank0[150]} = 32'h0;
    {bank3[151], bank2[151], bank1[151], bank0[151]} = 32'h0;
    {bank3[152], bank2[152], bank1[152], bank0[152]} = 32'h0;
    {bank3[153], bank2[153], bank1[153], bank0[153]} = 32'h0;
    {bank3[154], bank2[154], bank1[154], bank0[154]} = 32'h0;
    {bank3[155], bank2[155], bank1[155], bank0[155]} = 32'h0;
    {bank3[156], bank2[156], bank1[156], bank0[156]} = 32'h0;
    {bank3[157], bank2[157], bank1[157], bank0[157]} = 32'h0;
    {bank3[158], bank2[158], bank1[158], bank0[158]} = 32'h0;
    {bank3[159], bank2[159], bank1[159], bank0[159]} = 32'h0;
    {bank3[160], bank2[160], bank1[160], bank0[160]} = 32'h0;
    {bank3[161], bank2[161], bank1[161], bank0[161]} = 32'h0;
    {bank3[162], bank2[162], bank1[162], bank0[162]} = 32'h0;
    {bank3[163], bank2[163], bank1[163], bank0[163]} = 32'h0;
    {bank3[164], bank2[164], bank1[164], bank0[164]} = 32'h0;
    {bank3[165], bank2[165], bank1[165], bank0[165]} = 32'h0;
    {bank3[166], bank2[166], bank1[166], bank0[166]} = 32'h0;
    {bank3[167], bank2[167], bank1[167], bank0[167]} = 32'h0;
    {bank3[168], bank2[168], bank1[168], bank0[168]} = 32'h0;
    {bank3[169], bank2[169], bank1[169], bank0[169]} = 32'h0;
    {bank3[170], bank2[170], bank1[170], bank0[170]} = 32'h0;
    {bank3[171], bank2[171], bank1[171], bank0[171]} = 32'h0;
    {bank3[172], bank2[172], bank1[172], bank0[172]} = 32'h0;
    {bank3[173], bank2[173], bank1[173], bank0[173]} = 32'h0;
    {bank3[174], bank2[174], bank1[174], bank0[174]} = 32'h0;
    {bank3[175], bank2[175], bank1[175], bank0[175]} = 32'h0;
    {bank3[176], bank2[176], bank1[176], bank0[176]} = 32'h0;
    {bank3[177], bank2[177], bank1[177], bank0[177]} = 32'h0;
    {bank3[178], bank2[178], bank1[178], bank0[178]} = 32'h0;
    {bank3[179], bank2[179], bank1[179], bank0[179]} = 32'h0;
    {bank3[180], bank2[180], bank1[180], bank0[180]} = 32'h0;
    {bank3[181], bank2[181], bank1[181], bank0[181]} = 32'h0;
    {bank3[182], bank2[182], bank1[182], bank0[182]} = 32'h0;
    {bank3[183], bank2[183], bank1[183], bank0[183]} = 32'h0;
    {bank3[184], bank2[184], bank1[184], bank0[184]} = 32'h0;
    {bank3[185], bank2[185], bank1[185], bank0[185]} = 32'h0;
    {bank3[186], bank2[186], bank1[186], bank0[186]} = 32'h0;
    {bank3[187], bank2[187], bank1[187], bank0[187]} = 32'h0;
    {bank3[188], bank2[188], bank1[188], bank0[188]} = 32'h0;
    {bank3[189], bank2[189], bank1[189], bank0[189]} = 32'h0;
    {bank3[190], bank2[190], bank1[190], bank0[190]} = 32'h0;
    {bank3[191], bank2[191], bank1[191], bank0[191]} = 32'h0;
    {bank3[192], bank2[192], bank1[192], bank0[192]} = 32'h0;
    {bank3[193], bank2[193], bank1[193], bank0[193]} = 32'h0;
    {bank3[194], bank2[194], bank1[194], bank0[194]} = 32'h0;
    {bank3[195], bank2[195], bank1[195], bank0[195]} = 32'h0;
    {bank3[196], bank2[196], bank1[196], bank0[196]} = 32'h0;
    {bank3[197], bank2[197], bank1[197], bank0[197]} = 32'h0;
    {bank3[198], bank2[198], bank1[198], bank0[198]} = 32'h0;
    {bank3[199], bank2[199], bank1[199], bank0[199]} = 32'h0;
    {bank3[200], bank2[200], bank1[200], bank0[200]} = 32'h0;
    {bank3[201], bank2[201], bank1[201], bank0[201]} = 32'h0;
    {bank3[202], bank2[202], bank1[202], bank0[202]} = 32'h0;
    {bank3[203], bank2[203], bank1[203], bank0[203]} = 32'h0;
    {bank3[204], bank2[204], bank1[204], bank0[204]} = 32'h0;
    {bank3[205], bank2[205], bank1[205], bank0[205]} = 32'h0;
    {bank3[206], bank2[206], bank1[206], bank0[206]} = 32'h0;
    {bank3[207], bank2[207], bank1[207], bank0[207]} = 32'h0;
    {bank3[208], bank2[208], bank1[208], bank0[208]} = 32'h0;
    {bank3[209], bank2[209], bank1[209], bank0[209]} = 32'h0;
    {bank3[210], bank2[210], bank1[210], bank0[210]} = 32'h0;
    {bank3[211], bank2[211], bank1[211], bank0[211]} = 32'h0;
    {bank3[212], bank2[212], bank1[212], bank0[212]} = 32'h0;
    {bank3[213], bank2[213], bank1[213], bank0[213]} = 32'h0;
    {bank3[214], bank2[214], bank1[214], bank0[214]} = 32'h0;
    {bank3[215], bank2[215], bank1[215], bank0[215]} = 32'h0;
    {bank3[216], bank2[216], bank1[216], bank0[216]} = 32'h0;
    {bank3[217], bank2[217], bank1[217], bank0[217]} = 32'h0;
    {bank3[218], bank2[218], bank1[218], bank0[218]} = 32'h0;
    {bank3[219], bank2[219], bank1[219], bank0[219]} = 32'h0;
    {bank3[220], bank2[220], bank1[220], bank0[220]} = 32'h0;
    {bank3[221], bank2[221], bank1[221], bank0[221]} = 32'h0;
    {bank3[222], bank2[222], bank1[222], bank0[222]} = 32'h0;
    {bank3[223], bank2[223], bank1[223], bank0[223]} = 32'h0;
    {bank3[224], bank2[224], bank1[224], bank0[224]} = 32'h0;
    {bank3[225], bank2[225], bank1[225], bank0[225]} = 32'h0;
    {bank3[226], bank2[226], bank1[226], bank0[226]} = 32'h0;
    {bank3[227], bank2[227], bank1[227], bank0[227]} = 32'h0;
    {bank3[228], bank2[228], bank1[228], bank0[228]} = 32'h0;
    {bank3[229], bank2[229], bank1[229], bank0[229]} = 32'h0;
    {bank3[230], bank2[230], bank1[230], bank0[230]} = 32'h0;
    {bank3[231], bank2[231], bank1[231], bank0[231]} = 32'h0;
    {bank3[232], bank2[232], bank1[232], bank0[232]} = 32'h0;
    {bank3[233], bank2[233], bank1[233], bank0[233]} = 32'h0;
    {bank3[234], bank2[234], bank1[234], bank0[234]} = 32'h0;
    {bank3[235], bank2[235], bank1[235], bank0[235]} = 32'h0;
    {bank3[236], bank2[236], bank1[236], bank0[236]} = 32'h0;
    {bank3[237], bank2[237], bank1[237], bank0[237]} = 32'h0;
    {bank3[238], bank2[238], bank1[238], bank0[238]} = 32'h0;
    {bank3[239], bank2[239], bank1[239], bank0[239]} = 32'h0;
    {bank3[240], bank2[240], bank1[240], bank0[240]} = 32'h0;
    {bank3[241], bank2[241], bank1[241], bank0[241]} = 32'h0;
    {bank3[242], bank2[242], bank1[242], bank0[242]} = 32'h0;
    {bank3[243], bank2[243], bank1[243], bank0[243]} = 32'h0;
    {bank3[244], bank2[244], bank1[244], bank0[244]} = 32'h0;
    {bank3[245], bank2[245], bank1[245], bank0[245]} = 32'h0;
    {bank3[246], bank2[246], bank1[246], bank0[246]} = 32'h0;
    {bank3[247], bank2[247], bank1[247], bank0[247]} = 32'h0;
    {bank3[248], bank2[248], bank1[248], bank0[248]} = 32'h0;
    {bank3[249], bank2[249], bank1[249], bank0[249]} = 32'h0;
    {bank3[250], bank2[250], bank1[250], bank0[250]} = 32'h0;
    {bank3[251], bank2[251], bank1[251], bank0[251]} = 32'h0;
    {bank3[252], bank2[252], bank1[252], bank0[252]} = 32'h0;
    {bank3[253], bank2[253], bank1[253], bank0[253]} = 32'h0;
    {bank3[254], bank2[254], bank1[254], bank0[254]} = 32'h0;
    {bank3[255], bank2[255], bank1[255], bank0[255]} = 32'h0;
    {bank3[256], bank2[256], bank1[256], bank0[256]} = 32'h0;
    {bank3[257], bank2[257], bank1[257], bank0[257]} = 32'h0;
    {bank3[258], bank2[258], bank1[258], bank0[258]} = 32'h0;
    {bank3[259], bank2[259], bank1[259], bank0[259]} = 32'h0;
    {bank3[260], bank2[260], bank1[260], bank0[260]} = 32'h0;
    {bank3[261], bank2[261], bank1[261], bank0[261]} = 32'h0;
    {bank3[262], bank2[262], bank1[262], bank0[262]} = 32'h0;
    {bank3[263], bank2[263], bank1[263], bank0[263]} = 32'h0;
    {bank3[264], bank2[264], bank1[264], bank0[264]} = 32'h0;
    {bank3[265], bank2[265], bank1[265], bank0[265]} = 32'h0;
    {bank3[266], bank2[266], bank1[266], bank0[266]} = 32'h0;
    {bank3[267], bank2[267], bank1[267], bank0[267]} = 32'h0;
    {bank3[268], bank2[268], bank1[268], bank0[268]} = 32'h0;
    {bank3[269], bank2[269], bank1[269], bank0[269]} = 32'h0;
    {bank3[270], bank2[270], bank1[270], bank0[270]} = 32'h0;
    {bank3[271], bank2[271], bank1[271], bank0[271]} = 32'h0;
    {bank3[272], bank2[272], bank1[272], bank0[272]} = 32'h0;
    {bank3[273], bank2[273], bank1[273], bank0[273]} = 32'h0;
    {bank3[274], bank2[274], bank1[274], bank0[274]} = 32'h0;
    {bank3[275], bank2[275], bank1[275], bank0[275]} = 32'h0;
    {bank3[276], bank2[276], bank1[276], bank0[276]} = 32'h0;
    {bank3[277], bank2[277], bank1[277], bank0[277]} = 32'h0;
    {bank3[278], bank2[278], bank1[278], bank0[278]} = 32'h0;
    {bank3[279], bank2[279], bank1[279], bank0[279]} = 32'h0;
    {bank3[280], bank2[280], bank1[280], bank0[280]} = 32'h0;
    {bank3[281], bank2[281], bank1[281], bank0[281]} = 32'h0;
    {bank3[282], bank2[282], bank1[282], bank0[282]} = 32'h0;
    {bank3[283], bank2[283], bank1[283], bank0[283]} = 32'h0;
    {bank3[284], bank2[284], bank1[284], bank0[284]} = 32'h0;
    {bank3[285], bank2[285], bank1[285], bank0[285]} = 32'h0;
    {bank3[286], bank2[286], bank1[286], bank0[286]} = 32'h0;
    {bank3[287], bank2[287], bank1[287], bank0[287]} = 32'h0;
    {bank3[288], bank2[288], bank1[288], bank0[288]} = 32'h0;
    {bank3[289], bank2[289], bank1[289], bank0[289]} = 32'h0;
    {bank3[290], bank2[290], bank1[290], bank0[290]} = 32'h0;
    {bank3[291], bank2[291], bank1[291], bank0[291]} = 32'h0;
    {bank3[292], bank2[292], bank1[292], bank0[292]} = 32'h0;
    {bank3[293], bank2[293], bank1[293], bank0[293]} = 32'h0;
    {bank3[294], bank2[294], bank1[294], bank0[294]} = 32'h0;
    {bank3[295], bank2[295], bank1[295], bank0[295]} = 32'h0;
    {bank3[296], bank2[296], bank1[296], bank0[296]} = 32'h0;
    {bank3[297], bank2[297], bank1[297], bank0[297]} = 32'h0;
    {bank3[298], bank2[298], bank1[298], bank0[298]} = 32'h0;
    {bank3[299], bank2[299], bank1[299], bank0[299]} = 32'h0;
    {bank3[300], bank2[300], bank1[300], bank0[300]} = 32'h0;
    {bank3[301], bank2[301], bank1[301], bank0[301]} = 32'h0;
    {bank3[302], bank2[302], bank1[302], bank0[302]} = 32'h0;
    {bank3[303], bank2[303], bank1[303], bank0[303]} = 32'h0;
    {bank3[304], bank2[304], bank1[304], bank0[304]} = 32'h0;
    {bank3[305], bank2[305], bank1[305], bank0[305]} = 32'h0;
    {bank3[306], bank2[306], bank1[306], bank0[306]} = 32'h0;
    {bank3[307], bank2[307], bank1[307], bank0[307]} = 32'h0;
    {bank3[308], bank2[308], bank1[308], bank0[308]} = 32'h0;
    {bank3[309], bank2[309], bank1[309], bank0[309]} = 32'h0;
    {bank3[310], bank2[310], bank1[310], bank0[310]} = 32'h0;
    {bank3[311], bank2[311], bank1[311], bank0[311]} = 32'h0;
    {bank3[312], bank2[312], bank1[312], bank0[312]} = 32'h0;
    {bank3[313], bank2[313], bank1[313], bank0[313]} = 32'h0;
    {bank3[314], bank2[314], bank1[314], bank0[314]} = 32'h0;
    {bank3[315], bank2[315], bank1[315], bank0[315]} = 32'h0;
    {bank3[316], bank2[316], bank1[316], bank0[316]} = 32'h0;
    {bank3[317], bank2[317], bank1[317], bank0[317]} = 32'h0;
    {bank3[318], bank2[318], bank1[318], bank0[318]} = 32'h0;
    {bank3[319], bank2[319], bank1[319], bank0[319]} = 32'h0;
    {bank3[320], bank2[320], bank1[320], bank0[320]} = 32'h0;
    {bank3[321], bank2[321], bank1[321], bank0[321]} = 32'h0;
    {bank3[322], bank2[322], bank1[322], bank0[322]} = 32'h0;
    {bank3[323], bank2[323], bank1[323], bank0[323]} = 32'h0;
    {bank3[324], bank2[324], bank1[324], bank0[324]} = 32'h0;
    {bank3[325], bank2[325], bank1[325], bank0[325]} = 32'h0;
    {bank3[326], bank2[326], bank1[326], bank0[326]} = 32'h0;
    {bank3[327], bank2[327], bank1[327], bank0[327]} = 32'h0;
    {bank3[328], bank2[328], bank1[328], bank0[328]} = 32'h0;
    {bank3[329], bank2[329], bank1[329], bank0[329]} = 32'h0;
    {bank3[330], bank2[330], bank1[330], bank0[330]} = 32'h0;
    {bank3[331], bank2[331], bank1[331], bank0[331]} = 32'h0;
    {bank3[332], bank2[332], bank1[332], bank0[332]} = 32'h0;
    {bank3[333], bank2[333], bank1[333], bank0[333]} = 32'h0;
    {bank3[334], bank2[334], bank1[334], bank0[334]} = 32'h0;
    {bank3[335], bank2[335], bank1[335], bank0[335]} = 32'h0;
    {bank3[336], bank2[336], bank1[336], bank0[336]} = 32'h0;
    {bank3[337], bank2[337], bank1[337], bank0[337]} = 32'h0;
    {bank3[338], bank2[338], bank1[338], bank0[338]} = 32'h0;
    {bank3[339], bank2[339], bank1[339], bank0[339]} = 32'h0;
    {bank3[340], bank2[340], bank1[340], bank0[340]} = 32'h0;
    {bank3[341], bank2[341], bank1[341], bank0[341]} = 32'h0;
    {bank3[342], bank2[342], bank1[342], bank0[342]} = 32'h0;
    {bank3[343], bank2[343], bank1[343], bank0[343]} = 32'h0;
    {bank3[344], bank2[344], bank1[344], bank0[344]} = 32'h0;
    {bank3[345], bank2[345], bank1[345], bank0[345]} = 32'h0;
    {bank3[346], bank2[346], bank1[346], bank0[346]} = 32'h0;
    {bank3[347], bank2[347], bank1[347], bank0[347]} = 32'h0;
    {bank3[348], bank2[348], bank1[348], bank0[348]} = 32'h0;
    {bank3[349], bank2[349], bank1[349], bank0[349]} = 32'h0;
    {bank3[350], bank2[350], bank1[350], bank0[350]} = 32'h0;
    {bank3[351], bank2[351], bank1[351], bank0[351]} = 32'h0;
    {bank3[352], bank2[352], bank1[352], bank0[352]} = 32'h0;
    {bank3[353], bank2[353], bank1[353], bank0[353]} = 32'h0;
    {bank3[354], bank2[354], bank1[354], bank0[354]} = 32'h0;
    {bank3[355], bank2[355], bank1[355], bank0[355]} = 32'h0;
    {bank3[356], bank2[356], bank1[356], bank0[356]} = 32'h0;
    {bank3[357], bank2[357], bank1[357], bank0[357]} = 32'h0;
    {bank3[358], bank2[358], bank1[358], bank0[358]} = 32'h0;
    {bank3[359], bank2[359], bank1[359], bank0[359]} = 32'h0;
    {bank3[360], bank2[360], bank1[360], bank0[360]} = 32'h0;
    {bank3[361], bank2[361], bank1[361], bank0[361]} = 32'h0;
    {bank3[362], bank2[362], bank1[362], bank0[362]} = 32'h0;
    {bank3[363], bank2[363], bank1[363], bank0[363]} = 32'h0;
    {bank3[364], bank2[364], bank1[364], bank0[364]} = 32'h0;
    {bank3[365], bank2[365], bank1[365], bank0[365]} = 32'h0;
    {bank3[366], bank2[366], bank1[366], bank0[366]} = 32'h0;
    {bank3[367], bank2[367], bank1[367], bank0[367]} = 32'h0;
    {bank3[368], bank2[368], bank1[368], bank0[368]} = 32'h0;
    {bank3[369], bank2[369], bank1[369], bank0[369]} = 32'h0;
    {bank3[370], bank2[370], bank1[370], bank0[370]} = 32'h0;
    {bank3[371], bank2[371], bank1[371], bank0[371]} = 32'h0;
    {bank3[372], bank2[372], bank1[372], bank0[372]} = 32'h0;
    {bank3[373], bank2[373], bank1[373], bank0[373]} = 32'h0;
    {bank3[374], bank2[374], bank1[374], bank0[374]} = 32'h0;
    {bank3[375], bank2[375], bank1[375], bank0[375]} = 32'h0;
    {bank3[376], bank2[376], bank1[376], bank0[376]} = 32'h0;
    {bank3[377], bank2[377], bank1[377], bank0[377]} = 32'h0;
    {bank3[378], bank2[378], bank1[378], bank0[378]} = 32'h0;
    {bank3[379], bank2[379], bank1[379], bank0[379]} = 32'h0;
    {bank3[380], bank2[380], bank1[380], bank0[380]} = 32'h0;
    {bank3[381], bank2[381], bank1[381], bank0[381]} = 32'h0;
    {bank3[382], bank2[382], bank1[382], bank0[382]} = 32'h0;
    {bank3[383], bank2[383], bank1[383], bank0[383]} = 32'h0;
    {bank3[384], bank2[384], bank1[384], bank0[384]} = 32'h0;
    {bank3[385], bank2[385], bank1[385], bank0[385]} = 32'h0;
    {bank3[386], bank2[386], bank1[386], bank0[386]} = 32'h0;
    {bank3[387], bank2[387], bank1[387], bank0[387]} = 32'h0;
    {bank3[388], bank2[388], bank1[388], bank0[388]} = 32'h0;
    {bank3[389], bank2[389], bank1[389], bank0[389]} = 32'h0;
    {bank3[390], bank2[390], bank1[390], bank0[390]} = 32'h0;
    {bank3[391], bank2[391], bank1[391], bank0[391]} = 32'h0;
    {bank3[392], bank2[392], bank1[392], bank0[392]} = 32'h0;
    {bank3[393], bank2[393], bank1[393], bank0[393]} = 32'h0;
    {bank3[394], bank2[394], bank1[394], bank0[394]} = 32'h0;
    {bank3[395], bank2[395], bank1[395], bank0[395]} = 32'h0;
    {bank3[396], bank2[396], bank1[396], bank0[396]} = 32'h0;
    {bank3[397], bank2[397], bank1[397], bank0[397]} = 32'h0;
    {bank3[398], bank2[398], bank1[398], bank0[398]} = 32'h0;
    {bank3[399], bank2[399], bank1[399], bank0[399]} = 32'h0;
    {bank3[400], bank2[400], bank1[400], bank0[400]} = 32'h0;
    {bank3[401], bank2[401], bank1[401], bank0[401]} = 32'h0;
    {bank3[402], bank2[402], bank1[402], bank0[402]} = 32'h0;
    {bank3[403], bank2[403], bank1[403], bank0[403]} = 32'h0;
    {bank3[404], bank2[404], bank1[404], bank0[404]} = 32'h0;
    {bank3[405], bank2[405], bank1[405], bank0[405]} = 32'h0;
    {bank3[406], bank2[406], bank1[406], bank0[406]} = 32'h0;
    {bank3[407], bank2[407], bank1[407], bank0[407]} = 32'h0;
    {bank3[408], bank2[408], bank1[408], bank0[408]} = 32'h0;
    {bank3[409], bank2[409], bank1[409], bank0[409]} = 32'h0;
    {bank3[410], bank2[410], bank1[410], bank0[410]} = 32'h0;
    {bank3[411], bank2[411], bank1[411], bank0[411]} = 32'h0;
    {bank3[412], bank2[412], bank1[412], bank0[412]} = 32'h0;
    {bank3[413], bank2[413], bank1[413], bank0[413]} = 32'h0;
    {bank3[414], bank2[414], bank1[414], bank0[414]} = 32'h0;
    {bank3[415], bank2[415], bank1[415], bank0[415]} = 32'h0;
    {bank3[416], bank2[416], bank1[416], bank0[416]} = 32'h0;
    {bank3[417], bank2[417], bank1[417], bank0[417]} = 32'h0;
    {bank3[418], bank2[418], bank1[418], bank0[418]} = 32'h0;
    {bank3[419], bank2[419], bank1[419], bank0[419]} = 32'h0;
    {bank3[420], bank2[420], bank1[420], bank0[420]} = 32'h0;
    {bank3[421], bank2[421], bank1[421], bank0[421]} = 32'h0;
    {bank3[422], bank2[422], bank1[422], bank0[422]} = 32'h0;
    {bank3[423], bank2[423], bank1[423], bank0[423]} = 32'h0;
    {bank3[424], bank2[424], bank1[424], bank0[424]} = 32'h0;
    {bank3[425], bank2[425], bank1[425], bank0[425]} = 32'h0;
    {bank3[426], bank2[426], bank1[426], bank0[426]} = 32'h0;
    {bank3[427], bank2[427], bank1[427], bank0[427]} = 32'h0;
    {bank3[428], bank2[428], bank1[428], bank0[428]} = 32'h0;
    {bank3[429], bank2[429], bank1[429], bank0[429]} = 32'h0;
    {bank3[430], bank2[430], bank1[430], bank0[430]} = 32'h0;
    {bank3[431], bank2[431], bank1[431], bank0[431]} = 32'h0;
    {bank3[432], bank2[432], bank1[432], bank0[432]} = 32'h0;
    {bank3[433], bank2[433], bank1[433], bank0[433]} = 32'h0;
    {bank3[434], bank2[434], bank1[434], bank0[434]} = 32'h0;
    {bank3[435], bank2[435], bank1[435], bank0[435]} = 32'h0;
    {bank3[436], bank2[436], bank1[436], bank0[436]} = 32'h0;
    {bank3[437], bank2[437], bank1[437], bank0[437]} = 32'h0;
    {bank3[438], bank2[438], bank1[438], bank0[438]} = 32'h0;
    {bank3[439], bank2[439], bank1[439], bank0[439]} = 32'h0;
    {bank3[440], bank2[440], bank1[440], bank0[440]} = 32'h0;
    {bank3[441], bank2[441], bank1[441], bank0[441]} = 32'h0;
    {bank3[442], bank2[442], bank1[442], bank0[442]} = 32'h0;
    {bank3[443], bank2[443], bank1[443], bank0[443]} = 32'h0;
    {bank3[444], bank2[444], bank1[444], bank0[444]} = 32'h0;
    {bank3[445], bank2[445], bank1[445], bank0[445]} = 32'h0;
    {bank3[446], bank2[446], bank1[446], bank0[446]} = 32'h0;
    {bank3[447], bank2[447], bank1[447], bank0[447]} = 32'h0;
    {bank3[448], bank2[448], bank1[448], bank0[448]} = 32'h0;
    {bank3[449], bank2[449], bank1[449], bank0[449]} = 32'h0;
    {bank3[450], bank2[450], bank1[450], bank0[450]} = 32'h0;
    {bank3[451], bank2[451], bank1[451], bank0[451]} = 32'h0;
    {bank3[452], bank2[452], bank1[452], bank0[452]} = 32'h0;
    {bank3[453], bank2[453], bank1[453], bank0[453]} = 32'h0;
    {bank3[454], bank2[454], bank1[454], bank0[454]} = 32'h0;
    {bank3[455], bank2[455], bank1[455], bank0[455]} = 32'h0;
    {bank3[456], bank2[456], bank1[456], bank0[456]} = 32'h0;
    {bank3[457], bank2[457], bank1[457], bank0[457]} = 32'h0;
    {bank3[458], bank2[458], bank1[458], bank0[458]} = 32'h0;
    {bank3[459], bank2[459], bank1[459], bank0[459]} = 32'h0;
    {bank3[460], bank2[460], bank1[460], bank0[460]} = 32'h0;
    {bank3[461], bank2[461], bank1[461], bank0[461]} = 32'h0;
    {bank3[462], bank2[462], bank1[462], bank0[462]} = 32'h0;
    {bank3[463], bank2[463], bank1[463], bank0[463]} = 32'h0;
    {bank3[464], bank2[464], bank1[464], bank0[464]} = 32'h0;
    {bank3[465], bank2[465], bank1[465], bank0[465]} = 32'h0;
    {bank3[466], bank2[466], bank1[466], bank0[466]} = 32'h0;
    {bank3[467], bank2[467], bank1[467], bank0[467]} = 32'h0;
    {bank3[468], bank2[468], bank1[468], bank0[468]} = 32'h0;
    {bank3[469], bank2[469], bank1[469], bank0[469]} = 32'h0;
    {bank3[470], bank2[470], bank1[470], bank0[470]} = 32'h0;
    {bank3[471], bank2[471], bank1[471], bank0[471]} = 32'h0;
    {bank3[472], bank2[472], bank1[472], bank0[472]} = 32'h0;
    {bank3[473], bank2[473], bank1[473], bank0[473]} = 32'h0;
    {bank3[474], bank2[474], bank1[474], bank0[474]} = 32'h0;
    {bank3[475], bank2[475], bank1[475], bank0[475]} = 32'h0;
    {bank3[476], bank2[476], bank1[476], bank0[476]} = 32'h0;
    {bank3[477], bank2[477], bank1[477], bank0[477]} = 32'h0;
    {bank3[478], bank2[478], bank1[478], bank0[478]} = 32'h0;
    {bank3[479], bank2[479], bank1[479], bank0[479]} = 32'h0;
    {bank3[480], bank2[480], bank1[480], bank0[480]} = 32'h0;
    {bank3[481], bank2[481], bank1[481], bank0[481]} = 32'h0;
    {bank3[482], bank2[482], bank1[482], bank0[482]} = 32'h0;
    {bank3[483], bank2[483], bank1[483], bank0[483]} = 32'h0;
    {bank3[484], bank2[484], bank1[484], bank0[484]} = 32'h0;
    {bank3[485], bank2[485], bank1[485], bank0[485]} = 32'h0;
    {bank3[486], bank2[486], bank1[486], bank0[486]} = 32'h0;
    {bank3[487], bank2[487], bank1[487], bank0[487]} = 32'h0;
    {bank3[488], bank2[488], bank1[488], bank0[488]} = 32'h0;
    {bank3[489], bank2[489], bank1[489], bank0[489]} = 32'h0;
    {bank3[490], bank2[490], bank1[490], bank0[490]} = 32'h0;
    {bank3[491], bank2[491], bank1[491], bank0[491]} = 32'h0;
    {bank3[492], bank2[492], bank1[492], bank0[492]} = 32'h0;
    {bank3[493], bank2[493], bank1[493], bank0[493]} = 32'h0;
    {bank3[494], bank2[494], bank1[494], bank0[494]} = 32'h0;
    {bank3[495], bank2[495], bank1[495], bank0[495]} = 32'h0;
    {bank3[496], bank2[496], bank1[496], bank0[496]} = 32'h0;
    {bank3[497], bank2[497], bank1[497], bank0[497]} = 32'h0;
    {bank3[498], bank2[498], bank1[498], bank0[498]} = 32'h0;
    {bank3[499], bank2[499], bank1[499], bank0[499]} = 32'h0;
    {bank3[500], bank2[500], bank1[500], bank0[500]} = 32'h0;
    {bank3[501], bank2[501], bank1[501], bank0[501]} = 32'h0;
    {bank3[502], bank2[502], bank1[502], bank0[502]} = 32'h0;
    {bank3[503], bank2[503], bank1[503], bank0[503]} = 32'h0;
    {bank3[504], bank2[504], bank1[504], bank0[504]} = 32'h0;
    {bank3[505], bank2[505], bank1[505], bank0[505]} = 32'h0;
    {bank3[506], bank2[506], bank1[506], bank0[506]} = 32'h0;
    {bank3[507], bank2[507], bank1[507], bank0[507]} = 32'h0;
    {bank3[508], bank2[508], bank1[508], bank0[508]} = 32'h0;
    {bank3[509], bank2[509], bank1[509], bank0[509]} = 32'h0;
    {bank3[510], bank2[510], bank1[510], bank0[510]} = 32'h0;
    {bank3[511], bank2[511], bank1[511], bank0[511]} = 32'h0;
    {bank3[512], bank2[512], bank1[512], bank0[512]} = 32'h0;
    {bank3[513], bank2[513], bank1[513], bank0[513]} = 32'h0;
    {bank3[514], bank2[514], bank1[514], bank0[514]} = 32'h0;
    {bank3[515], bank2[515], bank1[515], bank0[515]} = 32'h0;
    {bank3[516], bank2[516], bank1[516], bank0[516]} = 32'h0;
    {bank3[517], bank2[517], bank1[517], bank0[517]} = 32'h0;
    {bank3[518], bank2[518], bank1[518], bank0[518]} = 32'h0;
    {bank3[519], bank2[519], bank1[519], bank0[519]} = 32'h0;
    {bank3[520], bank2[520], bank1[520], bank0[520]} = 32'h0;
    {bank3[521], bank2[521], bank1[521], bank0[521]} = 32'h0;
    {bank3[522], bank2[522], bank1[522], bank0[522]} = 32'h0;
    {bank3[523], bank2[523], bank1[523], bank0[523]} = 32'h0;
    {bank3[524], bank2[524], bank1[524], bank0[524]} = 32'h0;
    {bank3[525], bank2[525], bank1[525], bank0[525]} = 32'h0;
    {bank3[526], bank2[526], bank1[526], bank0[526]} = 32'h0;
    {bank3[527], bank2[527], bank1[527], bank0[527]} = 32'h0;
    {bank3[528], bank2[528], bank1[528], bank0[528]} = 32'h0;
    {bank3[529], bank2[529], bank1[529], bank0[529]} = 32'h0;
    {bank3[530], bank2[530], bank1[530], bank0[530]} = 32'h0;
    {bank3[531], bank2[531], bank1[531], bank0[531]} = 32'h0;
    {bank3[532], bank2[532], bank1[532], bank0[532]} = 32'h0;
    {bank3[533], bank2[533], bank1[533], bank0[533]} = 32'h0;
    {bank3[534], bank2[534], bank1[534], bank0[534]} = 32'h0;
    {bank3[535], bank2[535], bank1[535], bank0[535]} = 32'h0;
    {bank3[536], bank2[536], bank1[536], bank0[536]} = 32'h0;
    {bank3[537], bank2[537], bank1[537], bank0[537]} = 32'h0;
    {bank3[538], bank2[538], bank1[538], bank0[538]} = 32'h0;
    {bank3[539], bank2[539], bank1[539], bank0[539]} = 32'h0;
    {bank3[540], bank2[540], bank1[540], bank0[540]} = 32'h0;
    {bank3[541], bank2[541], bank1[541], bank0[541]} = 32'h0;
    {bank3[542], bank2[542], bank1[542], bank0[542]} = 32'h0;
    {bank3[543], bank2[543], bank1[543], bank0[543]} = 32'h0;
    {bank3[544], bank2[544], bank1[544], bank0[544]} = 32'h0;
    {bank3[545], bank2[545], bank1[545], bank0[545]} = 32'h0;
    {bank3[546], bank2[546], bank1[546], bank0[546]} = 32'h0;
    {bank3[547], bank2[547], bank1[547], bank0[547]} = 32'h0;
    {bank3[548], bank2[548], bank1[548], bank0[548]} = 32'h0;
    {bank3[549], bank2[549], bank1[549], bank0[549]} = 32'h0;
    {bank3[550], bank2[550], bank1[550], bank0[550]} = 32'h0;
    {bank3[551], bank2[551], bank1[551], bank0[551]} = 32'h0;
    {bank3[552], bank2[552], bank1[552], bank0[552]} = 32'h0;
    {bank3[553], bank2[553], bank1[553], bank0[553]} = 32'h0;
    {bank3[554], bank2[554], bank1[554], bank0[554]} = 32'h0;
    {bank3[555], bank2[555], bank1[555], bank0[555]} = 32'h0;
    {bank3[556], bank2[556], bank1[556], bank0[556]} = 32'h0;
    {bank3[557], bank2[557], bank1[557], bank0[557]} = 32'h0;
    {bank3[558], bank2[558], bank1[558], bank0[558]} = 32'h0;
    {bank3[559], bank2[559], bank1[559], bank0[559]} = 32'h0;
    {bank3[560], bank2[560], bank1[560], bank0[560]} = 32'h0;
    {bank3[561], bank2[561], bank1[561], bank0[561]} = 32'h0;
    {bank3[562], bank2[562], bank1[562], bank0[562]} = 32'h0;
    {bank3[563], bank2[563], bank1[563], bank0[563]} = 32'h0;
    {bank3[564], bank2[564], bank1[564], bank0[564]} = 32'h0;
    {bank3[565], bank2[565], bank1[565], bank0[565]} = 32'h0;
    {bank3[566], bank2[566], bank1[566], bank0[566]} = 32'h0;
    {bank3[567], bank2[567], bank1[567], bank0[567]} = 32'h0;
    {bank3[568], bank2[568], bank1[568], bank0[568]} = 32'h0;
    {bank3[569], bank2[569], bank1[569], bank0[569]} = 32'h0;
    {bank3[570], bank2[570], bank1[570], bank0[570]} = 32'h0;
    {bank3[571], bank2[571], bank1[571], bank0[571]} = 32'h0;
    {bank3[572], bank2[572], bank1[572], bank0[572]} = 32'h0;
    {bank3[573], bank2[573], bank1[573], bank0[573]} = 32'h0;
    {bank3[574], bank2[574], bank1[574], bank0[574]} = 32'h0;
    {bank3[575], bank2[575], bank1[575], bank0[575]} = 32'h0;
    {bank3[576], bank2[576], bank1[576], bank0[576]} = 32'h0;
    {bank3[577], bank2[577], bank1[577], bank0[577]} = 32'h0;
    {bank3[578], bank2[578], bank1[578], bank0[578]} = 32'h0;
    {bank3[579], bank2[579], bank1[579], bank0[579]} = 32'h0;
    {bank3[580], bank2[580], bank1[580], bank0[580]} = 32'h0;
    {bank3[581], bank2[581], bank1[581], bank0[581]} = 32'h0;
    {bank3[582], bank2[582], bank1[582], bank0[582]} = 32'h0;
    {bank3[583], bank2[583], bank1[583], bank0[583]} = 32'h0;
    {bank3[584], bank2[584], bank1[584], bank0[584]} = 32'h0;
    {bank3[585], bank2[585], bank1[585], bank0[585]} = 32'h0;
    {bank3[586], bank2[586], bank1[586], bank0[586]} = 32'h0;
    {bank3[587], bank2[587], bank1[587], bank0[587]} = 32'h0;
    {bank3[588], bank2[588], bank1[588], bank0[588]} = 32'h0;
    {bank3[589], bank2[589], bank1[589], bank0[589]} = 32'h0;
    {bank3[590], bank2[590], bank1[590], bank0[590]} = 32'h0;
    {bank3[591], bank2[591], bank1[591], bank0[591]} = 32'h0;
    {bank3[592], bank2[592], bank1[592], bank0[592]} = 32'h0;
    {bank3[593], bank2[593], bank1[593], bank0[593]} = 32'h0;
    {bank3[594], bank2[594], bank1[594], bank0[594]} = 32'h0;
    {bank3[595], bank2[595], bank1[595], bank0[595]} = 32'h0;
    {bank3[596], bank2[596], bank1[596], bank0[596]} = 32'h0;
    {bank3[597], bank2[597], bank1[597], bank0[597]} = 32'h0;
    {bank3[598], bank2[598], bank1[598], bank0[598]} = 32'h0;
    {bank3[599], bank2[599], bank1[599], bank0[599]} = 32'h0;
    {bank3[600], bank2[600], bank1[600], bank0[600]} = 32'h0;
    {bank3[601], bank2[601], bank1[601], bank0[601]} = 32'h0;
    {bank3[602], bank2[602], bank1[602], bank0[602]} = 32'h0;
    {bank3[603], bank2[603], bank1[603], bank0[603]} = 32'h0;
    {bank3[604], bank2[604], bank1[604], bank0[604]} = 32'h0;
    {bank3[605], bank2[605], bank1[605], bank0[605]} = 32'h0;
    {bank3[606], bank2[606], bank1[606], bank0[606]} = 32'h0;
    {bank3[607], bank2[607], bank1[607], bank0[607]} = 32'h0;
    {bank3[608], bank2[608], bank1[608], bank0[608]} = 32'h0;
    {bank3[609], bank2[609], bank1[609], bank0[609]} = 32'h0;
    {bank3[610], bank2[610], bank1[610], bank0[610]} = 32'h0;
    {bank3[611], bank2[611], bank1[611], bank0[611]} = 32'h0;
    {bank3[612], bank2[612], bank1[612], bank0[612]} = 32'h0;
    {bank3[613], bank2[613], bank1[613], bank0[613]} = 32'h0;
    {bank3[614], bank2[614], bank1[614], bank0[614]} = 32'h0;
    {bank3[615], bank2[615], bank1[615], bank0[615]} = 32'h0;
    {bank3[616], bank2[616], bank1[616], bank0[616]} = 32'h0;
    {bank3[617], bank2[617], bank1[617], bank0[617]} = 32'h0;
    {bank3[618], bank2[618], bank1[618], bank0[618]} = 32'h0;
    {bank3[619], bank2[619], bank1[619], bank0[619]} = 32'h0;
    {bank3[620], bank2[620], bank1[620], bank0[620]} = 32'h0;
    {bank3[621], bank2[621], bank1[621], bank0[621]} = 32'h0;
    {bank3[622], bank2[622], bank1[622], bank0[622]} = 32'h0;
    {bank3[623], bank2[623], bank1[623], bank0[623]} = 32'h0;
    {bank3[624], bank2[624], bank1[624], bank0[624]} = 32'h0;
    {bank3[625], bank2[625], bank1[625], bank0[625]} = 32'h0;
    {bank3[626], bank2[626], bank1[626], bank0[626]} = 32'h0;
    {bank3[627], bank2[627], bank1[627], bank0[627]} = 32'h0;
    {bank3[628], bank2[628], bank1[628], bank0[628]} = 32'h0;
    {bank3[629], bank2[629], bank1[629], bank0[629]} = 32'h0;
    {bank3[630], bank2[630], bank1[630], bank0[630]} = 32'h0;
    {bank3[631], bank2[631], bank1[631], bank0[631]} = 32'h0;
    {bank3[632], bank2[632], bank1[632], bank0[632]} = 32'h0;
    {bank3[633], bank2[633], bank1[633], bank0[633]} = 32'h0;
    {bank3[634], bank2[634], bank1[634], bank0[634]} = 32'h0;
    {bank3[635], bank2[635], bank1[635], bank0[635]} = 32'h0;
    {bank3[636], bank2[636], bank1[636], bank0[636]} = 32'h0;
    {bank3[637], bank2[637], bank1[637], bank0[637]} = 32'h0;
    {bank3[638], bank2[638], bank1[638], bank0[638]} = 32'h0;
    {bank3[639], bank2[639], bank1[639], bank0[639]} = 32'h0;
    {bank3[640], bank2[640], bank1[640], bank0[640]} = 32'h0;
    {bank3[641], bank2[641], bank1[641], bank0[641]} = 32'h0;
    {bank3[642], bank2[642], bank1[642], bank0[642]} = 32'h0;
    {bank3[643], bank2[643], bank1[643], bank0[643]} = 32'h0;
    {bank3[644], bank2[644], bank1[644], bank0[644]} = 32'h0;
    {bank3[645], bank2[645], bank1[645], bank0[645]} = 32'h0;
    {bank3[646], bank2[646], bank1[646], bank0[646]} = 32'h0;
    {bank3[647], bank2[647], bank1[647], bank0[647]} = 32'h0;
    {bank3[648], bank2[648], bank1[648], bank0[648]} = 32'h0;
    {bank3[649], bank2[649], bank1[649], bank0[649]} = 32'h0;
    {bank3[650], bank2[650], bank1[650], bank0[650]} = 32'h0;
    {bank3[651], bank2[651], bank1[651], bank0[651]} = 32'h0;
    {bank3[652], bank2[652], bank1[652], bank0[652]} = 32'h0;
    {bank3[653], bank2[653], bank1[653], bank0[653]} = 32'h0;
    {bank3[654], bank2[654], bank1[654], bank0[654]} = 32'h0;
    {bank3[655], bank2[655], bank1[655], bank0[655]} = 32'h0;
    {bank3[656], bank2[656], bank1[656], bank0[656]} = 32'h0;
    {bank3[657], bank2[657], bank1[657], bank0[657]} = 32'h0;
    {bank3[658], bank2[658], bank1[658], bank0[658]} = 32'h0;
    {bank3[659], bank2[659], bank1[659], bank0[659]} = 32'h0;
    {bank3[660], bank2[660], bank1[660], bank0[660]} = 32'h0;
    {bank3[661], bank2[661], bank1[661], bank0[661]} = 32'h0;
    {bank3[662], bank2[662], bank1[662], bank0[662]} = 32'h0;
    {bank3[663], bank2[663], bank1[663], bank0[663]} = 32'h0;
    {bank3[664], bank2[664], bank1[664], bank0[664]} = 32'h0;
    {bank3[665], bank2[665], bank1[665], bank0[665]} = 32'h0;
    {bank3[666], bank2[666], bank1[666], bank0[666]} = 32'h0;
    {bank3[667], bank2[667], bank1[667], bank0[667]} = 32'h0;
    {bank3[668], bank2[668], bank1[668], bank0[668]} = 32'h0;
    {bank3[669], bank2[669], bank1[669], bank0[669]} = 32'h0;
    {bank3[670], bank2[670], bank1[670], bank0[670]} = 32'h0;
    {bank3[671], bank2[671], bank1[671], bank0[671]} = 32'h0;
    {bank3[672], bank2[672], bank1[672], bank0[672]} = 32'h0;
    {bank3[673], bank2[673], bank1[673], bank0[673]} = 32'h0;
    {bank3[674], bank2[674], bank1[674], bank0[674]} = 32'h0;
    {bank3[675], bank2[675], bank1[675], bank0[675]} = 32'h0;
    {bank3[676], bank2[676], bank1[676], bank0[676]} = 32'h0;
    {bank3[677], bank2[677], bank1[677], bank0[677]} = 32'h0;
    {bank3[678], bank2[678], bank1[678], bank0[678]} = 32'h0;
    {bank3[679], bank2[679], bank1[679], bank0[679]} = 32'h0;
    {bank3[680], bank2[680], bank1[680], bank0[680]} = 32'h0;
    {bank3[681], bank2[681], bank1[681], bank0[681]} = 32'h0;
    {bank3[682], bank2[682], bank1[682], bank0[682]} = 32'h0;
    {bank3[683], bank2[683], bank1[683], bank0[683]} = 32'h0;
    {bank3[684], bank2[684], bank1[684], bank0[684]} = 32'h0;
    {bank3[685], bank2[685], bank1[685], bank0[685]} = 32'h0;
    {bank3[686], bank2[686], bank1[686], bank0[686]} = 32'h0;
    {bank3[687], bank2[687], bank1[687], bank0[687]} = 32'h0;
    {bank3[688], bank2[688], bank1[688], bank0[688]} = 32'h0;
    {bank3[689], bank2[689], bank1[689], bank0[689]} = 32'h0;
    {bank3[690], bank2[690], bank1[690], bank0[690]} = 32'h0;
    {bank3[691], bank2[691], bank1[691], bank0[691]} = 32'h0;
    {bank3[692], bank2[692], bank1[692], bank0[692]} = 32'h0;
    {bank3[693], bank2[693], bank1[693], bank0[693]} = 32'h0;
    {bank3[694], bank2[694], bank1[694], bank0[694]} = 32'h0;
    {bank3[695], bank2[695], bank1[695], bank0[695]} = 32'h0;
    {bank3[696], bank2[696], bank1[696], bank0[696]} = 32'h0;
    {bank3[697], bank2[697], bank1[697], bank0[697]} = 32'h0;
    {bank3[698], bank2[698], bank1[698], bank0[698]} = 32'h0;
    {bank3[699], bank2[699], bank1[699], bank0[699]} = 32'h0;
    {bank3[700], bank2[700], bank1[700], bank0[700]} = 32'h0;
    {bank3[701], bank2[701], bank1[701], bank0[701]} = 32'h0;
    {bank3[702], bank2[702], bank1[702], bank0[702]} = 32'h0;
    {bank3[703], bank2[703], bank1[703], bank0[703]} = 32'h0;
    {bank3[704], bank2[704], bank1[704], bank0[704]} = 32'h0;
    {bank3[705], bank2[705], bank1[705], bank0[705]} = 32'h0;
    {bank3[706], bank2[706], bank1[706], bank0[706]} = 32'h0;
    {bank3[707], bank2[707], bank1[707], bank0[707]} = 32'h0;
    {bank3[708], bank2[708], bank1[708], bank0[708]} = 32'h0;
    {bank3[709], bank2[709], bank1[709], bank0[709]} = 32'h0;
    {bank3[710], bank2[710], bank1[710], bank0[710]} = 32'h0;
    {bank3[711], bank2[711], bank1[711], bank0[711]} = 32'h0;
    {bank3[712], bank2[712], bank1[712], bank0[712]} = 32'h0;
    {bank3[713], bank2[713], bank1[713], bank0[713]} = 32'h0;
    {bank3[714], bank2[714], bank1[714], bank0[714]} = 32'h0;
    {bank3[715], bank2[715], bank1[715], bank0[715]} = 32'h0;
    {bank3[716], bank2[716], bank1[716], bank0[716]} = 32'h0;
    {bank3[717], bank2[717], bank1[717], bank0[717]} = 32'h0;
    {bank3[718], bank2[718], bank1[718], bank0[718]} = 32'h0;
    {bank3[719], bank2[719], bank1[719], bank0[719]} = 32'h0;
    {bank3[720], bank2[720], bank1[720], bank0[720]} = 32'h0;
    {bank3[721], bank2[721], bank1[721], bank0[721]} = 32'h0;
    {bank3[722], bank2[722], bank1[722], bank0[722]} = 32'h0;
    {bank3[723], bank2[723], bank1[723], bank0[723]} = 32'h0;
    {bank3[724], bank2[724], bank1[724], bank0[724]} = 32'h0;
    {bank3[725], bank2[725], bank1[725], bank0[725]} = 32'h0;
    {bank3[726], bank2[726], bank1[726], bank0[726]} = 32'h0;
    {bank3[727], bank2[727], bank1[727], bank0[727]} = 32'h0;
    {bank3[728], bank2[728], bank1[728], bank0[728]} = 32'h0;
    {bank3[729], bank2[729], bank1[729], bank0[729]} = 32'h0;
    {bank3[730], bank2[730], bank1[730], bank0[730]} = 32'h0;
    {bank3[731], bank2[731], bank1[731], bank0[731]} = 32'h0;
    {bank3[732], bank2[732], bank1[732], bank0[732]} = 32'h0;
    {bank3[733], bank2[733], bank1[733], bank0[733]} = 32'h0;
    {bank3[734], bank2[734], bank1[734], bank0[734]} = 32'h0;
    {bank3[735], bank2[735], bank1[735], bank0[735]} = 32'h0;
    {bank3[736], bank2[736], bank1[736], bank0[736]} = 32'h0;
    {bank3[737], bank2[737], bank1[737], bank0[737]} = 32'h0;
    {bank3[738], bank2[738], bank1[738], bank0[738]} = 32'h0;
    {bank3[739], bank2[739], bank1[739], bank0[739]} = 32'h0;
    {bank3[740], bank2[740], bank1[740], bank0[740]} = 32'h0;
    {bank3[741], bank2[741], bank1[741], bank0[741]} = 32'h0;
    {bank3[742], bank2[742], bank1[742], bank0[742]} = 32'h0;
    {bank3[743], bank2[743], bank1[743], bank0[743]} = 32'h0;
    {bank3[744], bank2[744], bank1[744], bank0[744]} = 32'h0;
    {bank3[745], bank2[745], bank1[745], bank0[745]} = 32'h0;
    {bank3[746], bank2[746], bank1[746], bank0[746]} = 32'h0;
    {bank3[747], bank2[747], bank1[747], bank0[747]} = 32'h0;
    {bank3[748], bank2[748], bank1[748], bank0[748]} = 32'h0;
    {bank3[749], bank2[749], bank1[749], bank0[749]} = 32'h0;
    {bank3[750], bank2[750], bank1[750], bank0[750]} = 32'h0;
    {bank3[751], bank2[751], bank1[751], bank0[751]} = 32'h0;
    {bank3[752], bank2[752], bank1[752], bank0[752]} = 32'h0;
    {bank3[753], bank2[753], bank1[753], bank0[753]} = 32'h0;
    {bank3[754], bank2[754], bank1[754], bank0[754]} = 32'h0;
    {bank3[755], bank2[755], bank1[755], bank0[755]} = 32'h0;
    {bank3[756], bank2[756], bank1[756], bank0[756]} = 32'h0;
    {bank3[757], bank2[757], bank1[757], bank0[757]} = 32'h0;
    {bank3[758], bank2[758], bank1[758], bank0[758]} = 32'h0;
    {bank3[759], bank2[759], bank1[759], bank0[759]} = 32'h0;
    {bank3[760], bank2[760], bank1[760], bank0[760]} = 32'h0;
    {bank3[761], bank2[761], bank1[761], bank0[761]} = 32'h0;
    {bank3[762], bank2[762], bank1[762], bank0[762]} = 32'h0;
    {bank3[763], bank2[763], bank1[763], bank0[763]} = 32'h0;
    {bank3[764], bank2[764], bank1[764], bank0[764]} = 32'h0;
    {bank3[765], bank2[765], bank1[765], bank0[765]} = 32'h0;
    {bank3[766], bank2[766], bank1[766], bank0[766]} = 32'h0;
    {bank3[767], bank2[767], bank1[767], bank0[767]} = 32'h0;
    {bank3[768], bank2[768], bank1[768], bank0[768]} = 32'h0;
    {bank3[769], bank2[769], bank1[769], bank0[769]} = 32'h0;
    {bank3[770], bank2[770], bank1[770], bank0[770]} = 32'h0;
    {bank3[771], bank2[771], bank1[771], bank0[771]} = 32'h0;
    {bank3[772], bank2[772], bank1[772], bank0[772]} = 32'h0;
    {bank3[773], bank2[773], bank1[773], bank0[773]} = 32'h0;
    {bank3[774], bank2[774], bank1[774], bank0[774]} = 32'h0;
    {bank3[775], bank2[775], bank1[775], bank0[775]} = 32'h0;
    {bank3[776], bank2[776], bank1[776], bank0[776]} = 32'h0;
    {bank3[777], bank2[777], bank1[777], bank0[777]} = 32'h0;
    {bank3[778], bank2[778], bank1[778], bank0[778]} = 32'h0;
    {bank3[779], bank2[779], bank1[779], bank0[779]} = 32'h0;
    {bank3[780], bank2[780], bank1[780], bank0[780]} = 32'h0;
    {bank3[781], bank2[781], bank1[781], bank0[781]} = 32'h0;
    {bank3[782], bank2[782], bank1[782], bank0[782]} = 32'h0;
    {bank3[783], bank2[783], bank1[783], bank0[783]} = 32'h0;
    {bank3[784], bank2[784], bank1[784], bank0[784]} = 32'h0;
    {bank3[785], bank2[785], bank1[785], bank0[785]} = 32'h0;
    {bank3[786], bank2[786], bank1[786], bank0[786]} = 32'h0;
    {bank3[787], bank2[787], bank1[787], bank0[787]} = 32'h0;
    {bank3[788], bank2[788], bank1[788], bank0[788]} = 32'h0;
    {bank3[789], bank2[789], bank1[789], bank0[789]} = 32'h0;
    {bank3[790], bank2[790], bank1[790], bank0[790]} = 32'h0;
    {bank3[791], bank2[791], bank1[791], bank0[791]} = 32'h0;
    {bank3[792], bank2[792], bank1[792], bank0[792]} = 32'h0;
    {bank3[793], bank2[793], bank1[793], bank0[793]} = 32'h0;
    {bank3[794], bank2[794], bank1[794], bank0[794]} = 32'h0;
    {bank3[795], bank2[795], bank1[795], bank0[795]} = 32'h0;
    {bank3[796], bank2[796], bank1[796], bank0[796]} = 32'h0;
    {bank3[797], bank2[797], bank1[797], bank0[797]} = 32'h0;
    {bank3[798], bank2[798], bank1[798], bank0[798]} = 32'h0;
    {bank3[799], bank2[799], bank1[799], bank0[799]} = 32'h0;
    {bank3[800], bank2[800], bank1[800], bank0[800]} = 32'h0;
    {bank3[801], bank2[801], bank1[801], bank0[801]} = 32'h0;
    {bank3[802], bank2[802], bank1[802], bank0[802]} = 32'h0;
    {bank3[803], bank2[803], bank1[803], bank0[803]} = 32'h0;
    {bank3[804], bank2[804], bank1[804], bank0[804]} = 32'h0;
    {bank3[805], bank2[805], bank1[805], bank0[805]} = 32'h0;
    {bank3[806], bank2[806], bank1[806], bank0[806]} = 32'h0;
    {bank3[807], bank2[807], bank1[807], bank0[807]} = 32'h0;
    {bank3[808], bank2[808], bank1[808], bank0[808]} = 32'h0;
    {bank3[809], bank2[809], bank1[809], bank0[809]} = 32'h0;
    {bank3[810], bank2[810], bank1[810], bank0[810]} = 32'h0;
    {bank3[811], bank2[811], bank1[811], bank0[811]} = 32'h0;
    {bank3[812], bank2[812], bank1[812], bank0[812]} = 32'h0;
    {bank3[813], bank2[813], bank1[813], bank0[813]} = 32'h0;
    {bank3[814], bank2[814], bank1[814], bank0[814]} = 32'h0;
    {bank3[815], bank2[815], bank1[815], bank0[815]} = 32'h0;
    {bank3[816], bank2[816], bank1[816], bank0[816]} = 32'h0;
    {bank3[817], bank2[817], bank1[817], bank0[817]} = 32'h0;
    {bank3[818], bank2[818], bank1[818], bank0[818]} = 32'h0;
    {bank3[819], bank2[819], bank1[819], bank0[819]} = 32'h0;
    {bank3[820], bank2[820], bank1[820], bank0[820]} = 32'h0;
    {bank3[821], bank2[821], bank1[821], bank0[821]} = 32'h0;
    {bank3[822], bank2[822], bank1[822], bank0[822]} = 32'h0;
    {bank3[823], bank2[823], bank1[823], bank0[823]} = 32'h0;
    {bank3[824], bank2[824], bank1[824], bank0[824]} = 32'h0;
    {bank3[825], bank2[825], bank1[825], bank0[825]} = 32'h0;
    {bank3[826], bank2[826], bank1[826], bank0[826]} = 32'h0;
    {bank3[827], bank2[827], bank1[827], bank0[827]} = 32'h0;
    {bank3[828], bank2[828], bank1[828], bank0[828]} = 32'h0;
    {bank3[829], bank2[829], bank1[829], bank0[829]} = 32'h0;
    {bank3[830], bank2[830], bank1[830], bank0[830]} = 32'h0;
    {bank3[831], bank2[831], bank1[831], bank0[831]} = 32'h0;
    {bank3[832], bank2[832], bank1[832], bank0[832]} = 32'h0;
    {bank3[833], bank2[833], bank1[833], bank0[833]} = 32'h0;
    {bank3[834], bank2[834], bank1[834], bank0[834]} = 32'h0;
    {bank3[835], bank2[835], bank1[835], bank0[835]} = 32'h0;
    {bank3[836], bank2[836], bank1[836], bank0[836]} = 32'h0;
    {bank3[837], bank2[837], bank1[837], bank0[837]} = 32'h0;
    {bank3[838], bank2[838], bank1[838], bank0[838]} = 32'h0;
    {bank3[839], bank2[839], bank1[839], bank0[839]} = 32'h0;
    {bank3[840], bank2[840], bank1[840], bank0[840]} = 32'h0;
    {bank3[841], bank2[841], bank1[841], bank0[841]} = 32'h0;
    {bank3[842], bank2[842], bank1[842], bank0[842]} = 32'h0;
    {bank3[843], bank2[843], bank1[843], bank0[843]} = 32'h0;
    {bank3[844], bank2[844], bank1[844], bank0[844]} = 32'h0;
    {bank3[845], bank2[845], bank1[845], bank0[845]} = 32'h0;
    {bank3[846], bank2[846], bank1[846], bank0[846]} = 32'h0;
    {bank3[847], bank2[847], bank1[847], bank0[847]} = 32'h0;
    {bank3[848], bank2[848], bank1[848], bank0[848]} = 32'h0;
    {bank3[849], bank2[849], bank1[849], bank0[849]} = 32'h0;
    {bank3[850], bank2[850], bank1[850], bank0[850]} = 32'h0;
    {bank3[851], bank2[851], bank1[851], bank0[851]} = 32'h0;
    {bank3[852], bank2[852], bank1[852], bank0[852]} = 32'h0;
    {bank3[853], bank2[853], bank1[853], bank0[853]} = 32'h0;
    {bank3[854], bank2[854], bank1[854], bank0[854]} = 32'h0;
    {bank3[855], bank2[855], bank1[855], bank0[855]} = 32'h0;
    {bank3[856], bank2[856], bank1[856], bank0[856]} = 32'h0;
    {bank3[857], bank2[857], bank1[857], bank0[857]} = 32'h0;
    {bank3[858], bank2[858], bank1[858], bank0[858]} = 32'h0;
    {bank3[859], bank2[859], bank1[859], bank0[859]} = 32'h0;
    {bank3[860], bank2[860], bank1[860], bank0[860]} = 32'h0;
    {bank3[861], bank2[861], bank1[861], bank0[861]} = 32'h0;
    {bank3[862], bank2[862], bank1[862], bank0[862]} = 32'h0;
    {bank3[863], bank2[863], bank1[863], bank0[863]} = 32'h0;
    {bank3[864], bank2[864], bank1[864], bank0[864]} = 32'h0;
    {bank3[865], bank2[865], bank1[865], bank0[865]} = 32'h0;
    {bank3[866], bank2[866], bank1[866], bank0[866]} = 32'h0;
    {bank3[867], bank2[867], bank1[867], bank0[867]} = 32'h0;
    {bank3[868], bank2[868], bank1[868], bank0[868]} = 32'h0;
    {bank3[869], bank2[869], bank1[869], bank0[869]} = 32'h0;
    {bank3[870], bank2[870], bank1[870], bank0[870]} = 32'h0;
    {bank3[871], bank2[871], bank1[871], bank0[871]} = 32'h0;
    {bank3[872], bank2[872], bank1[872], bank0[872]} = 32'h0;
    {bank3[873], bank2[873], bank1[873], bank0[873]} = 32'h0;
    {bank3[874], bank2[874], bank1[874], bank0[874]} = 32'h0;
    {bank3[875], bank2[875], bank1[875], bank0[875]} = 32'h0;
    {bank3[876], bank2[876], bank1[876], bank0[876]} = 32'h0;
    {bank3[877], bank2[877], bank1[877], bank0[877]} = 32'h0;
    {bank3[878], bank2[878], bank1[878], bank0[878]} = 32'h0;
    {bank3[879], bank2[879], bank1[879], bank0[879]} = 32'h0;
    {bank3[880], bank2[880], bank1[880], bank0[880]} = 32'h0;
    {bank3[881], bank2[881], bank1[881], bank0[881]} = 32'h0;
    {bank3[882], bank2[882], bank1[882], bank0[882]} = 32'h0;
    {bank3[883], bank2[883], bank1[883], bank0[883]} = 32'h0;
    {bank3[884], bank2[884], bank1[884], bank0[884]} = 32'h0;
    {bank3[885], bank2[885], bank1[885], bank0[885]} = 32'h0;
    {bank3[886], bank2[886], bank1[886], bank0[886]} = 32'h0;
    {bank3[887], bank2[887], bank1[887], bank0[887]} = 32'h0;
    {bank3[888], bank2[888], bank1[888], bank0[888]} = 32'h0;
    {bank3[889], bank2[889], bank1[889], bank0[889]} = 32'h0;
    {bank3[890], bank2[890], bank1[890], bank0[890]} = 32'h0;
    {bank3[891], bank2[891], bank1[891], bank0[891]} = 32'h0;
    {bank3[892], bank2[892], bank1[892], bank0[892]} = 32'h0;
    {bank3[893], bank2[893], bank1[893], bank0[893]} = 32'h0;
    {bank3[894], bank2[894], bank1[894], bank0[894]} = 32'h0;
    {bank3[895], bank2[895], bank1[895], bank0[895]} = 32'h0;
    {bank3[896], bank2[896], bank1[896], bank0[896]} = 32'h0;
    {bank3[897], bank2[897], bank1[897], bank0[897]} = 32'h0;
    {bank3[898], bank2[898], bank1[898], bank0[898]} = 32'h0;
    {bank3[899], bank2[899], bank1[899], bank0[899]} = 32'h0;
    {bank3[900], bank2[900], bank1[900], bank0[900]} = 32'h0;
    {bank3[901], bank2[901], bank1[901], bank0[901]} = 32'h0;
    {bank3[902], bank2[902], bank1[902], bank0[902]} = 32'h0;
    {bank3[903], bank2[903], bank1[903], bank0[903]} = 32'h0;
    {bank3[904], bank2[904], bank1[904], bank0[904]} = 32'h0;
    {bank3[905], bank2[905], bank1[905], bank0[905]} = 32'h0;
    {bank3[906], bank2[906], bank1[906], bank0[906]} = 32'h0;
    {bank3[907], bank2[907], bank1[907], bank0[907]} = 32'h0;
    {bank3[908], bank2[908], bank1[908], bank0[908]} = 32'h0;
    {bank3[909], bank2[909], bank1[909], bank0[909]} = 32'h0;
    {bank3[910], bank2[910], bank1[910], bank0[910]} = 32'h0;
    {bank3[911], bank2[911], bank1[911], bank0[911]} = 32'h0;
    {bank3[912], bank2[912], bank1[912], bank0[912]} = 32'h0;
    {bank3[913], bank2[913], bank1[913], bank0[913]} = 32'h0;
    {bank3[914], bank2[914], bank1[914], bank0[914]} = 32'h0;
    {bank3[915], bank2[915], bank1[915], bank0[915]} = 32'h0;
    {bank3[916], bank2[916], bank1[916], bank0[916]} = 32'h0;
    {bank3[917], bank2[917], bank1[917], bank0[917]} = 32'h0;
    {bank3[918], bank2[918], bank1[918], bank0[918]} = 32'h0;
    {bank3[919], bank2[919], bank1[919], bank0[919]} = 32'h0;
    {bank3[920], bank2[920], bank1[920], bank0[920]} = 32'h0;
    {bank3[921], bank2[921], bank1[921], bank0[921]} = 32'h0;
    {bank3[922], bank2[922], bank1[922], bank0[922]} = 32'h0;
    {bank3[923], bank2[923], bank1[923], bank0[923]} = 32'h0;
    {bank3[924], bank2[924], bank1[924], bank0[924]} = 32'h0;
    {bank3[925], bank2[925], bank1[925], bank0[925]} = 32'h0;
    {bank3[926], bank2[926], bank1[926], bank0[926]} = 32'h0;
    {bank3[927], bank2[927], bank1[927], bank0[927]} = 32'h0;
    {bank3[928], bank2[928], bank1[928], bank0[928]} = 32'h0;
    {bank3[929], bank2[929], bank1[929], bank0[929]} = 32'h0;
    {bank3[930], bank2[930], bank1[930], bank0[930]} = 32'h0;
    {bank3[931], bank2[931], bank1[931], bank0[931]} = 32'h0;
    {bank3[932], bank2[932], bank1[932], bank0[932]} = 32'h0;
    {bank3[933], bank2[933], bank1[933], bank0[933]} = 32'h0;
    {bank3[934], bank2[934], bank1[934], bank0[934]} = 32'h0;
    {bank3[935], bank2[935], bank1[935], bank0[935]} = 32'h0;
    {bank3[936], bank2[936], bank1[936], bank0[936]} = 32'h0;
    {bank3[937], bank2[937], bank1[937], bank0[937]} = 32'h0;
    {bank3[938], bank2[938], bank1[938], bank0[938]} = 32'h0;
    {bank3[939], bank2[939], bank1[939], bank0[939]} = 32'h0;
    {bank3[940], bank2[940], bank1[940], bank0[940]} = 32'h0;
    {bank3[941], bank2[941], bank1[941], bank0[941]} = 32'h0;
    {bank3[942], bank2[942], bank1[942], bank0[942]} = 32'h0;
    {bank3[943], bank2[943], bank1[943], bank0[943]} = 32'h0;
    {bank3[944], bank2[944], bank1[944], bank0[944]} = 32'h0;
    {bank3[945], bank2[945], bank1[945], bank0[945]} = 32'h0;
    {bank3[946], bank2[946], bank1[946], bank0[946]} = 32'h0;
    {bank3[947], bank2[947], bank1[947], bank0[947]} = 32'h0;
    {bank3[948], bank2[948], bank1[948], bank0[948]} = 32'h0;
    {bank3[949], bank2[949], bank1[949], bank0[949]} = 32'h0;
    {bank3[950], bank2[950], bank1[950], bank0[950]} = 32'h0;
    {bank3[951], bank2[951], bank1[951], bank0[951]} = 32'h0;
    {bank3[952], bank2[952], bank1[952], bank0[952]} = 32'h0;
    {bank3[953], bank2[953], bank1[953], bank0[953]} = 32'h0;
    {bank3[954], bank2[954], bank1[954], bank0[954]} = 32'h0;
    {bank3[955], bank2[955], bank1[955], bank0[955]} = 32'h0;
    {bank3[956], bank2[956], bank1[956], bank0[956]} = 32'h0;
    {bank3[957], bank2[957], bank1[957], bank0[957]} = 32'h0;
    {bank3[958], bank2[958], bank1[958], bank0[958]} = 32'h0;
    {bank3[959], bank2[959], bank1[959], bank0[959]} = 32'h0;
    {bank3[960], bank2[960], bank1[960], bank0[960]} = 32'h0;
    {bank3[961], bank2[961], bank1[961], bank0[961]} = 32'h0;
    {bank3[962], bank2[962], bank1[962], bank0[962]} = 32'h0;
    {bank3[963], bank2[963], bank1[963], bank0[963]} = 32'h0;
    {bank3[964], bank2[964], bank1[964], bank0[964]} = 32'h0;
    {bank3[965], bank2[965], bank1[965], bank0[965]} = 32'h0;
    {bank3[966], bank2[966], bank1[966], bank0[966]} = 32'h0;
    {bank3[967], bank2[967], bank1[967], bank0[967]} = 32'h0;
    {bank3[968], bank2[968], bank1[968], bank0[968]} = 32'h0;
    {bank3[969], bank2[969], bank1[969], bank0[969]} = 32'h0;
    {bank3[970], bank2[970], bank1[970], bank0[970]} = 32'h0;
    {bank3[971], bank2[971], bank1[971], bank0[971]} = 32'h0;
    {bank3[972], bank2[972], bank1[972], bank0[972]} = 32'h0;
    {bank3[973], bank2[973], bank1[973], bank0[973]} = 32'h0;
    {bank3[974], bank2[974], bank1[974], bank0[974]} = 32'h0;
    {bank3[975], bank2[975], bank1[975], bank0[975]} = 32'h0;
    {bank3[976], bank2[976], bank1[976], bank0[976]} = 32'h0;
    {bank3[977], bank2[977], bank1[977], bank0[977]} = 32'h0;
    {bank3[978], bank2[978], bank1[978], bank0[978]} = 32'h0;
    {bank3[979], bank2[979], bank1[979], bank0[979]} = 32'h0;
    {bank3[980], bank2[980], bank1[980], bank0[980]} = 32'h0;
    {bank3[981], bank2[981], bank1[981], bank0[981]} = 32'h0;
    {bank3[982], bank2[982], bank1[982], bank0[982]} = 32'h0;
    {bank3[983], bank2[983], bank1[983], bank0[983]} = 32'h0;
    {bank3[984], bank2[984], bank1[984], bank0[984]} = 32'h0;
    {bank3[985], bank2[985], bank1[985], bank0[985]} = 32'h0;
    {bank3[986], bank2[986], bank1[986], bank0[986]} = 32'h0;
    {bank3[987], bank2[987], bank1[987], bank0[987]} = 32'h0;
    {bank3[988], bank2[988], bank1[988], bank0[988]} = 32'h0;
    {bank3[989], bank2[989], bank1[989], bank0[989]} = 32'h0;
    {bank3[990], bank2[990], bank1[990], bank0[990]} = 32'h0;
    {bank3[991], bank2[991], bank1[991], bank0[991]} = 32'h0;
    {bank3[992], bank2[992], bank1[992], bank0[992]} = 32'h0;
    {bank3[993], bank2[993], bank1[993], bank0[993]} = 32'h0;
    {bank3[994], bank2[994], bank1[994], bank0[994]} = 32'h0;
    {bank3[995], bank2[995], bank1[995], bank0[995]} = 32'h0;
    {bank3[996], bank2[996], bank1[996], bank0[996]} = 32'h0;
    {bank3[997], bank2[997], bank1[997], bank0[997]} = 32'h0;
    {bank3[998], bank2[998], bank1[998], bank0[998]} = 32'h0;
    {bank3[999], bank2[999], bank1[999], bank0[999]} = 32'h0;
    {bank3[1000], bank2[1000], bank1[1000], bank0[1000]} = 32'h0;
    {bank3[1001], bank2[1001], bank1[1001], bank0[1001]} = 32'h0;
    {bank3[1002], bank2[1002], bank1[1002], bank0[1002]} = 32'h0;
    {bank3[1003], bank2[1003], bank1[1003], bank0[1003]} = 32'h0;
    {bank3[1004], bank2[1004], bank1[1004], bank0[1004]} = 32'h0;
    {bank3[1005], bank2[1005], bank1[1005], bank0[1005]} = 32'h0;
    {bank3[1006], bank2[1006], bank1[1006], bank0[1006]} = 32'h0;
    {bank3[1007], bank2[1007], bank1[1007], bank0[1007]} = 32'h0;
    {bank3[1008], bank2[1008], bank1[1008], bank0[1008]} = 32'h0;
    {bank3[1009], bank2[1009], bank1[1009], bank0[1009]} = 32'h0;
    {bank3[1010], bank2[1010], bank1[1010], bank0[1010]} = 32'h0;
    {bank3[1011], bank2[1011], bank1[1011], bank0[1011]} = 32'h0;
    {bank3[1012], bank2[1012], bank1[1012], bank0[1012]} = 32'h0;
    {bank3[1013], bank2[1013], bank1[1013], bank0[1013]} = 32'h0;
    {bank3[1014], bank2[1014], bank1[1014], bank0[1014]} = 32'h0;
    {bank3[1015], bank2[1015], bank1[1015], bank0[1015]} = 32'h0;
    {bank3[1016], bank2[1016], bank1[1016], bank0[1016]} = 32'h0;
    {bank3[1017], bank2[1017], bank1[1017], bank0[1017]} = 32'h0;
    {bank3[1018], bank2[1018], bank1[1018], bank0[1018]} = 32'h0;
    {bank3[1019], bank2[1019], bank1[1019], bank0[1019]} = 32'h0;
    {bank3[1020], bank2[1020], bank1[1020], bank0[1020]} = 32'h0;
    {bank3[1021], bank2[1021], bank1[1021], bank0[1021]} = 32'h0;
    {bank3[1022], bank2[1022], bank1[1022], bank0[1022]} = 32'h0;
    {bank3[1023], bank2[1023], bank1[1023], bank0[1023]} = 32'h0;
    {bank3[1024], bank2[1024], bank1[1024], bank0[1024]} = 32'h0;
    {bank3[1025], bank2[1025], bank1[1025], bank0[1025]} = 32'h0;
    {bank3[1026], bank2[1026], bank1[1026], bank0[1026]} = 32'h0;
    {bank3[1027], bank2[1027], bank1[1027], bank0[1027]} = 32'h0;
    {bank3[1028], bank2[1028], bank1[1028], bank0[1028]} = 32'h0;
    {bank3[1029], bank2[1029], bank1[1029], bank0[1029]} = 32'h0;
    {bank3[1030], bank2[1030], bank1[1030], bank0[1030]} = 32'h0;
    {bank3[1031], bank2[1031], bank1[1031], bank0[1031]} = 32'h0;
    {bank3[1032], bank2[1032], bank1[1032], bank0[1032]} = 32'h0;
    {bank3[1033], bank2[1033], bank1[1033], bank0[1033]} = 32'h0;
    {bank3[1034], bank2[1034], bank1[1034], bank0[1034]} = 32'h0;
    {bank3[1035], bank2[1035], bank1[1035], bank0[1035]} = 32'h0;
    {bank3[1036], bank2[1036], bank1[1036], bank0[1036]} = 32'h0;
    {bank3[1037], bank2[1037], bank1[1037], bank0[1037]} = 32'h0;
    {bank3[1038], bank2[1038], bank1[1038], bank0[1038]} = 32'h0;
    {bank3[1039], bank2[1039], bank1[1039], bank0[1039]} = 32'h0;
    {bank3[1040], bank2[1040], bank1[1040], bank0[1040]} = 32'h0;
    {bank3[1041], bank2[1041], bank1[1041], bank0[1041]} = 32'h0;
    {bank3[1042], bank2[1042], bank1[1042], bank0[1042]} = 32'h0;
    {bank3[1043], bank2[1043], bank1[1043], bank0[1043]} = 32'h0;
    {bank3[1044], bank2[1044], bank1[1044], bank0[1044]} = 32'h0;
    {bank3[1045], bank2[1045], bank1[1045], bank0[1045]} = 32'h0;
    {bank3[1046], bank2[1046], bank1[1046], bank0[1046]} = 32'h0;
    {bank3[1047], bank2[1047], bank1[1047], bank0[1047]} = 32'h0;
    {bank3[1048], bank2[1048], bank1[1048], bank0[1048]} = 32'h0;
    {bank3[1049], bank2[1049], bank1[1049], bank0[1049]} = 32'h0;
    {bank3[1050], bank2[1050], bank1[1050], bank0[1050]} = 32'h0;
    {bank3[1051], bank2[1051], bank1[1051], bank0[1051]} = 32'h0;
    {bank3[1052], bank2[1052], bank1[1052], bank0[1052]} = 32'h0;
    {bank3[1053], bank2[1053], bank1[1053], bank0[1053]} = 32'h0;
    {bank3[1054], bank2[1054], bank1[1054], bank0[1054]} = 32'h0;
    {bank3[1055], bank2[1055], bank1[1055], bank0[1055]} = 32'h0;
    {bank3[1056], bank2[1056], bank1[1056], bank0[1056]} = 32'h0;
    {bank3[1057], bank2[1057], bank1[1057], bank0[1057]} = 32'h0;
    {bank3[1058], bank2[1058], bank1[1058], bank0[1058]} = 32'h0;
    {bank3[1059], bank2[1059], bank1[1059], bank0[1059]} = 32'h0;
    {bank3[1060], bank2[1060], bank1[1060], bank0[1060]} = 32'h0;
    {bank3[1061], bank2[1061], bank1[1061], bank0[1061]} = 32'h0;
    {bank3[1062], bank2[1062], bank1[1062], bank0[1062]} = 32'h0;
    {bank3[1063], bank2[1063], bank1[1063], bank0[1063]} = 32'h0;
    {bank3[1064], bank2[1064], bank1[1064], bank0[1064]} = 32'h0;
    {bank3[1065], bank2[1065], bank1[1065], bank0[1065]} = 32'h0;
    {bank3[1066], bank2[1066], bank1[1066], bank0[1066]} = 32'h0;
    {bank3[1067], bank2[1067], bank1[1067], bank0[1067]} = 32'h0;
    {bank3[1068], bank2[1068], bank1[1068], bank0[1068]} = 32'h0;
    {bank3[1069], bank2[1069], bank1[1069], bank0[1069]} = 32'h0;
    {bank3[1070], bank2[1070], bank1[1070], bank0[1070]} = 32'h0;
    {bank3[1071], bank2[1071], bank1[1071], bank0[1071]} = 32'h0;
    {bank3[1072], bank2[1072], bank1[1072], bank0[1072]} = 32'h0;
    {bank3[1073], bank2[1073], bank1[1073], bank0[1073]} = 32'h0;
    {bank3[1074], bank2[1074], bank1[1074], bank0[1074]} = 32'h0;
    {bank3[1075], bank2[1075], bank1[1075], bank0[1075]} = 32'h0;
    {bank3[1076], bank2[1076], bank1[1076], bank0[1076]} = 32'h0;
    {bank3[1077], bank2[1077], bank1[1077], bank0[1077]} = 32'h0;
    {bank3[1078], bank2[1078], bank1[1078], bank0[1078]} = 32'h0;
    {bank3[1079], bank2[1079], bank1[1079], bank0[1079]} = 32'h0;
    {bank3[1080], bank2[1080], bank1[1080], bank0[1080]} = 32'h0;
    {bank3[1081], bank2[1081], bank1[1081], bank0[1081]} = 32'h0;
    {bank3[1082], bank2[1082], bank1[1082], bank0[1082]} = 32'h0;
    {bank3[1083], bank2[1083], bank1[1083], bank0[1083]} = 32'h0;
    {bank3[1084], bank2[1084], bank1[1084], bank0[1084]} = 32'h0;
    {bank3[1085], bank2[1085], bank1[1085], bank0[1085]} = 32'h0;
    {bank3[1086], bank2[1086], bank1[1086], bank0[1086]} = 32'h0;
    {bank3[1087], bank2[1087], bank1[1087], bank0[1087]} = 32'h0;
    {bank3[1088], bank2[1088], bank1[1088], bank0[1088]} = 32'h0;
    {bank3[1089], bank2[1089], bank1[1089], bank0[1089]} = 32'h0;
    {bank3[1090], bank2[1090], bank1[1090], bank0[1090]} = 32'h0;
    {bank3[1091], bank2[1091], bank1[1091], bank0[1091]} = 32'h0;
    {bank3[1092], bank2[1092], bank1[1092], bank0[1092]} = 32'h0;
    {bank3[1093], bank2[1093], bank1[1093], bank0[1093]} = 32'h0;
    {bank3[1094], bank2[1094], bank1[1094], bank0[1094]} = 32'h0;
    {bank3[1095], bank2[1095], bank1[1095], bank0[1095]} = 32'h0;
    {bank3[1096], bank2[1096], bank1[1096], bank0[1096]} = 32'h0;
    {bank3[1097], bank2[1097], bank1[1097], bank0[1097]} = 32'h0;
    {bank3[1098], bank2[1098], bank1[1098], bank0[1098]} = 32'h0;
    {bank3[1099], bank2[1099], bank1[1099], bank0[1099]} = 32'h0;
    {bank3[1100], bank2[1100], bank1[1100], bank0[1100]} = 32'h0;
    {bank3[1101], bank2[1101], bank1[1101], bank0[1101]} = 32'h0;
    {bank3[1102], bank2[1102], bank1[1102], bank0[1102]} = 32'h0;
    {bank3[1103], bank2[1103], bank1[1103], bank0[1103]} = 32'h0;
    {bank3[1104], bank2[1104], bank1[1104], bank0[1104]} = 32'h0;
    {bank3[1105], bank2[1105], bank1[1105], bank0[1105]} = 32'h0;
    {bank3[1106], bank2[1106], bank1[1106], bank0[1106]} = 32'h0;
    {bank3[1107], bank2[1107], bank1[1107], bank0[1107]} = 32'h0;
    {bank3[1108], bank2[1108], bank1[1108], bank0[1108]} = 32'h0;
    {bank3[1109], bank2[1109], bank1[1109], bank0[1109]} = 32'h0;
    {bank3[1110], bank2[1110], bank1[1110], bank0[1110]} = 32'h0;
    {bank3[1111], bank2[1111], bank1[1111], bank0[1111]} = 32'h0;
    {bank3[1112], bank2[1112], bank1[1112], bank0[1112]} = 32'h0;
    {bank3[1113], bank2[1113], bank1[1113], bank0[1113]} = 32'h0;
    {bank3[1114], bank2[1114], bank1[1114], bank0[1114]} = 32'h0;
    {bank3[1115], bank2[1115], bank1[1115], bank0[1115]} = 32'h0;
    {bank3[1116], bank2[1116], bank1[1116], bank0[1116]} = 32'h0;
    {bank3[1117], bank2[1117], bank1[1117], bank0[1117]} = 32'h0;
    {bank3[1118], bank2[1118], bank1[1118], bank0[1118]} = 32'h0;
    {bank3[1119], bank2[1119], bank1[1119], bank0[1119]} = 32'h0;
    {bank3[1120], bank2[1120], bank1[1120], bank0[1120]} = 32'h0;
    {bank3[1121], bank2[1121], bank1[1121], bank0[1121]} = 32'h0;
    {bank3[1122], bank2[1122], bank1[1122], bank0[1122]} = 32'h0;
    {bank3[1123], bank2[1123], bank1[1123], bank0[1123]} = 32'h0;
    {bank3[1124], bank2[1124], bank1[1124], bank0[1124]} = 32'h0;
    {bank3[1125], bank2[1125], bank1[1125], bank0[1125]} = 32'h0;
    {bank3[1126], bank2[1126], bank1[1126], bank0[1126]} = 32'h0;
    {bank3[1127], bank2[1127], bank1[1127], bank0[1127]} = 32'h0;
    {bank3[1128], bank2[1128], bank1[1128], bank0[1128]} = 32'h0;
    {bank3[1129], bank2[1129], bank1[1129], bank0[1129]} = 32'h0;
    {bank3[1130], bank2[1130], bank1[1130], bank0[1130]} = 32'h0;
    {bank3[1131], bank2[1131], bank1[1131], bank0[1131]} = 32'h0;
    {bank3[1132], bank2[1132], bank1[1132], bank0[1132]} = 32'h0;
    {bank3[1133], bank2[1133], bank1[1133], bank0[1133]} = 32'h0;
    {bank3[1134], bank2[1134], bank1[1134], bank0[1134]} = 32'h0;
    {bank3[1135], bank2[1135], bank1[1135], bank0[1135]} = 32'h0;
    {bank3[1136], bank2[1136], bank1[1136], bank0[1136]} = 32'h0;
    {bank3[1137], bank2[1137], bank1[1137], bank0[1137]} = 32'h0;
    {bank3[1138], bank2[1138], bank1[1138], bank0[1138]} = 32'h0;
    {bank3[1139], bank2[1139], bank1[1139], bank0[1139]} = 32'h0;
    {bank3[1140], bank2[1140], bank1[1140], bank0[1140]} = 32'h0;
    {bank3[1141], bank2[1141], bank1[1141], bank0[1141]} = 32'h0;
    {bank3[1142], bank2[1142], bank1[1142], bank0[1142]} = 32'h0;
    {bank3[1143], bank2[1143], bank1[1143], bank0[1143]} = 32'h0;
    {bank3[1144], bank2[1144], bank1[1144], bank0[1144]} = 32'h0;
    {bank3[1145], bank2[1145], bank1[1145], bank0[1145]} = 32'h0;
    {bank3[1146], bank2[1146], bank1[1146], bank0[1146]} = 32'h0;
    {bank3[1147], bank2[1147], bank1[1147], bank0[1147]} = 32'h0;
    {bank3[1148], bank2[1148], bank1[1148], bank0[1148]} = 32'h0;
    {bank3[1149], bank2[1149], bank1[1149], bank0[1149]} = 32'h0;
    {bank3[1150], bank2[1150], bank1[1150], bank0[1150]} = 32'h0;
    {bank3[1151], bank2[1151], bank1[1151], bank0[1151]} = 32'h0;
    {bank3[1152], bank2[1152], bank1[1152], bank0[1152]} = 32'h0;
    {bank3[1153], bank2[1153], bank1[1153], bank0[1153]} = 32'h0;
    {bank3[1154], bank2[1154], bank1[1154], bank0[1154]} = 32'h0;
    {bank3[1155], bank2[1155], bank1[1155], bank0[1155]} = 32'h0;
    {bank3[1156], bank2[1156], bank1[1156], bank0[1156]} = 32'h0;
    {bank3[1157], bank2[1157], bank1[1157], bank0[1157]} = 32'h0;
    {bank3[1158], bank2[1158], bank1[1158], bank0[1158]} = 32'h0;
    {bank3[1159], bank2[1159], bank1[1159], bank0[1159]} = 32'h0;
    {bank3[1160], bank2[1160], bank1[1160], bank0[1160]} = 32'h0;
    {bank3[1161], bank2[1161], bank1[1161], bank0[1161]} = 32'h0;
    {bank3[1162], bank2[1162], bank1[1162], bank0[1162]} = 32'h0;
    {bank3[1163], bank2[1163], bank1[1163], bank0[1163]} = 32'h0;
    {bank3[1164], bank2[1164], bank1[1164], bank0[1164]} = 32'h0;
    {bank3[1165], bank2[1165], bank1[1165], bank0[1165]} = 32'h0;
    {bank3[1166], bank2[1166], bank1[1166], bank0[1166]} = 32'h0;
    {bank3[1167], bank2[1167], bank1[1167], bank0[1167]} = 32'h0;
    {bank3[1168], bank2[1168], bank1[1168], bank0[1168]} = 32'h0;
    {bank3[1169], bank2[1169], bank1[1169], bank0[1169]} = 32'h0;
    {bank3[1170], bank2[1170], bank1[1170], bank0[1170]} = 32'h0;
    {bank3[1171], bank2[1171], bank1[1171], bank0[1171]} = 32'h0;
    {bank3[1172], bank2[1172], bank1[1172], bank0[1172]} = 32'h0;
    {bank3[1173], bank2[1173], bank1[1173], bank0[1173]} = 32'h0;
    {bank3[1174], bank2[1174], bank1[1174], bank0[1174]} = 32'h0;
    {bank3[1175], bank2[1175], bank1[1175], bank0[1175]} = 32'h0;
    {bank3[1176], bank2[1176], bank1[1176], bank0[1176]} = 32'h0;
    {bank3[1177], bank2[1177], bank1[1177], bank0[1177]} = 32'h0;
    {bank3[1178], bank2[1178], bank1[1178], bank0[1178]} = 32'h0;
    {bank3[1179], bank2[1179], bank1[1179], bank0[1179]} = 32'h0;
    {bank3[1180], bank2[1180], bank1[1180], bank0[1180]} = 32'h0;
    {bank3[1181], bank2[1181], bank1[1181], bank0[1181]} = 32'h0;
    {bank3[1182], bank2[1182], bank1[1182], bank0[1182]} = 32'h0;
    {bank3[1183], bank2[1183], bank1[1183], bank0[1183]} = 32'h0;
    {bank3[1184], bank2[1184], bank1[1184], bank0[1184]} = 32'h0;
    {bank3[1185], bank2[1185], bank1[1185], bank0[1185]} = 32'h0;
    {bank3[1186], bank2[1186], bank1[1186], bank0[1186]} = 32'h0;
    {bank3[1187], bank2[1187], bank1[1187], bank0[1187]} = 32'h0;
    {bank3[1188], bank2[1188], bank1[1188], bank0[1188]} = 32'h0;
    {bank3[1189], bank2[1189], bank1[1189], bank0[1189]} = 32'h0;
    {bank3[1190], bank2[1190], bank1[1190], bank0[1190]} = 32'h0;
    {bank3[1191], bank2[1191], bank1[1191], bank0[1191]} = 32'h0;
    {bank3[1192], bank2[1192], bank1[1192], bank0[1192]} = 32'h0;
    {bank3[1193], bank2[1193], bank1[1193], bank0[1193]} = 32'h0;
    {bank3[1194], bank2[1194], bank1[1194], bank0[1194]} = 32'h0;
    {bank3[1195], bank2[1195], bank1[1195], bank0[1195]} = 32'h0;
    {bank3[1196], bank2[1196], bank1[1196], bank0[1196]} = 32'h0;
    {bank3[1197], bank2[1197], bank1[1197], bank0[1197]} = 32'h0;
    {bank3[1198], bank2[1198], bank1[1198], bank0[1198]} = 32'h0;
    {bank3[1199], bank2[1199], bank1[1199], bank0[1199]} = 32'h0;
    {bank3[1200], bank2[1200], bank1[1200], bank0[1200]} = 32'h0;
    {bank3[1201], bank2[1201], bank1[1201], bank0[1201]} = 32'h0;
    {bank3[1202], bank2[1202], bank1[1202], bank0[1202]} = 32'h0;
    {bank3[1203], bank2[1203], bank1[1203], bank0[1203]} = 32'h0;
    {bank3[1204], bank2[1204], bank1[1204], bank0[1204]} = 32'h0;
    {bank3[1205], bank2[1205], bank1[1205], bank0[1205]} = 32'h0;
    {bank3[1206], bank2[1206], bank1[1206], bank0[1206]} = 32'h0;
    {bank3[1207], bank2[1207], bank1[1207], bank0[1207]} = 32'h0;
    {bank3[1208], bank2[1208], bank1[1208], bank0[1208]} = 32'h0;
    {bank3[1209], bank2[1209], bank1[1209], bank0[1209]} = 32'h0;
    {bank3[1210], bank2[1210], bank1[1210], bank0[1210]} = 32'h0;
    {bank3[1211], bank2[1211], bank1[1211], bank0[1211]} = 32'h0;
    {bank3[1212], bank2[1212], bank1[1212], bank0[1212]} = 32'h0;
    {bank3[1213], bank2[1213], bank1[1213], bank0[1213]} = 32'h0;
    {bank3[1214], bank2[1214], bank1[1214], bank0[1214]} = 32'h0;
    {bank3[1215], bank2[1215], bank1[1215], bank0[1215]} = 32'h0;
    {bank3[1216], bank2[1216], bank1[1216], bank0[1216]} = 32'h0;
    {bank3[1217], bank2[1217], bank1[1217], bank0[1217]} = 32'h0;
    {bank3[1218], bank2[1218], bank1[1218], bank0[1218]} = 32'h0;
    {bank3[1219], bank2[1219], bank1[1219], bank0[1219]} = 32'h0;
    {bank3[1220], bank2[1220], bank1[1220], bank0[1220]} = 32'h0;
    {bank3[1221], bank2[1221], bank1[1221], bank0[1221]} = 32'h0;
    {bank3[1222], bank2[1222], bank1[1222], bank0[1222]} = 32'h0;
    {bank3[1223], bank2[1223], bank1[1223], bank0[1223]} = 32'h0;
    {bank3[1224], bank2[1224], bank1[1224], bank0[1224]} = 32'h0;
    {bank3[1225], bank2[1225], bank1[1225], bank0[1225]} = 32'h0;
    {bank3[1226], bank2[1226], bank1[1226], bank0[1226]} = 32'h0;
    {bank3[1227], bank2[1227], bank1[1227], bank0[1227]} = 32'h0;
    {bank3[1228], bank2[1228], bank1[1228], bank0[1228]} = 32'h0;
    {bank3[1229], bank2[1229], bank1[1229], bank0[1229]} = 32'h0;
    {bank3[1230], bank2[1230], bank1[1230], bank0[1230]} = 32'h0;
    {bank3[1231], bank2[1231], bank1[1231], bank0[1231]} = 32'h0;
    {bank3[1232], bank2[1232], bank1[1232], bank0[1232]} = 32'h0;
    {bank3[1233], bank2[1233], bank1[1233], bank0[1233]} = 32'h0;
    {bank3[1234], bank2[1234], bank1[1234], bank0[1234]} = 32'h0;
    {bank3[1235], bank2[1235], bank1[1235], bank0[1235]} = 32'h0;
    {bank3[1236], bank2[1236], bank1[1236], bank0[1236]} = 32'h0;
    {bank3[1237], bank2[1237], bank1[1237], bank0[1237]} = 32'h0;
    {bank3[1238], bank2[1238], bank1[1238], bank0[1238]} = 32'h0;
    {bank3[1239], bank2[1239], bank1[1239], bank0[1239]} = 32'h0;
    {bank3[1240], bank2[1240], bank1[1240], bank0[1240]} = 32'h0;
    {bank3[1241], bank2[1241], bank1[1241], bank0[1241]} = 32'h0;
    {bank3[1242], bank2[1242], bank1[1242], bank0[1242]} = 32'h0;
    {bank3[1243], bank2[1243], bank1[1243], bank0[1243]} = 32'h0;
    {bank3[1244], bank2[1244], bank1[1244], bank0[1244]} = 32'h0;
    {bank3[1245], bank2[1245], bank1[1245], bank0[1245]} = 32'h0;
    {bank3[1246], bank2[1246], bank1[1246], bank0[1246]} = 32'h0;
    {bank3[1247], bank2[1247], bank1[1247], bank0[1247]} = 32'h0;
    {bank3[1248], bank2[1248], bank1[1248], bank0[1248]} = 32'h0;
    {bank3[1249], bank2[1249], bank1[1249], bank0[1249]} = 32'h0;
    {bank3[1250], bank2[1250], bank1[1250], bank0[1250]} = 32'h0;
    {bank3[1251], bank2[1251], bank1[1251], bank0[1251]} = 32'h0;
    {bank3[1252], bank2[1252], bank1[1252], bank0[1252]} = 32'h0;
    {bank3[1253], bank2[1253], bank1[1253], bank0[1253]} = 32'h0;
    {bank3[1254], bank2[1254], bank1[1254], bank0[1254]} = 32'h0;
    {bank3[1255], bank2[1255], bank1[1255], bank0[1255]} = 32'h0;
    {bank3[1256], bank2[1256], bank1[1256], bank0[1256]} = 32'h0;
    {bank3[1257], bank2[1257], bank1[1257], bank0[1257]} = 32'h0;
    {bank3[1258], bank2[1258], bank1[1258], bank0[1258]} = 32'h0;
    {bank3[1259], bank2[1259], bank1[1259], bank0[1259]} = 32'h0;
    {bank3[1260], bank2[1260], bank1[1260], bank0[1260]} = 32'h0;
    {bank3[1261], bank2[1261], bank1[1261], bank0[1261]} = 32'h0;
    {bank3[1262], bank2[1262], bank1[1262], bank0[1262]} = 32'h0;
    {bank3[1263], bank2[1263], bank1[1263], bank0[1263]} = 32'h0;
    {bank3[1264], bank2[1264], bank1[1264], bank0[1264]} = 32'h0;
    {bank3[1265], bank2[1265], bank1[1265], bank0[1265]} = 32'h0;
    {bank3[1266], bank2[1266], bank1[1266], bank0[1266]} = 32'h0;
    {bank3[1267], bank2[1267], bank1[1267], bank0[1267]} = 32'h0;
    {bank3[1268], bank2[1268], bank1[1268], bank0[1268]} = 32'h0;
    {bank3[1269], bank2[1269], bank1[1269], bank0[1269]} = 32'h0;
    {bank3[1270], bank2[1270], bank1[1270], bank0[1270]} = 32'h0;
    {bank3[1271], bank2[1271], bank1[1271], bank0[1271]} = 32'h0;
    {bank3[1272], bank2[1272], bank1[1272], bank0[1272]} = 32'h0;
    {bank3[1273], bank2[1273], bank1[1273], bank0[1273]} = 32'h0;
    {bank3[1274], bank2[1274], bank1[1274], bank0[1274]} = 32'h0;
    {bank3[1275], bank2[1275], bank1[1275], bank0[1275]} = 32'h0;
    {bank3[1276], bank2[1276], bank1[1276], bank0[1276]} = 32'h0;
    {bank3[1277], bank2[1277], bank1[1277], bank0[1277]} = 32'h0;
    {bank3[1278], bank2[1278], bank1[1278], bank0[1278]} = 32'h0;
    {bank3[1279], bank2[1279], bank1[1279], bank0[1279]} = 32'h0;
    {bank3[1280], bank2[1280], bank1[1280], bank0[1280]} = 32'h0;
    {bank3[1281], bank2[1281], bank1[1281], bank0[1281]} = 32'h0;
    {bank3[1282], bank2[1282], bank1[1282], bank0[1282]} = 32'h0;
    {bank3[1283], bank2[1283], bank1[1283], bank0[1283]} = 32'h0;
    {bank3[1284], bank2[1284], bank1[1284], bank0[1284]} = 32'h0;
    {bank3[1285], bank2[1285], bank1[1285], bank0[1285]} = 32'h0;
    {bank3[1286], bank2[1286], bank1[1286], bank0[1286]} = 32'h0;
    {bank3[1287], bank2[1287], bank1[1287], bank0[1287]} = 32'h0;
    {bank3[1288], bank2[1288], bank1[1288], bank0[1288]} = 32'h0;
    {bank3[1289], bank2[1289], bank1[1289], bank0[1289]} = 32'h0;
    {bank3[1290], bank2[1290], bank1[1290], bank0[1290]} = 32'h0;
    {bank3[1291], bank2[1291], bank1[1291], bank0[1291]} = 32'h0;
    {bank3[1292], bank2[1292], bank1[1292], bank0[1292]} = 32'h0;
    {bank3[1293], bank2[1293], bank1[1293], bank0[1293]} = 32'h0;
    {bank3[1294], bank2[1294], bank1[1294], bank0[1294]} = 32'h0;
    {bank3[1295], bank2[1295], bank1[1295], bank0[1295]} = 32'h0;
    {bank3[1296], bank2[1296], bank1[1296], bank0[1296]} = 32'h0;
    {bank3[1297], bank2[1297], bank1[1297], bank0[1297]} = 32'h0;
    {bank3[1298], bank2[1298], bank1[1298], bank0[1298]} = 32'h0;
    {bank3[1299], bank2[1299], bank1[1299], bank0[1299]} = 32'h0;
    {bank3[1300], bank2[1300], bank1[1300], bank0[1300]} = 32'h0;
    {bank3[1301], bank2[1301], bank1[1301], bank0[1301]} = 32'h0;
    {bank3[1302], bank2[1302], bank1[1302], bank0[1302]} = 32'h0;
    {bank3[1303], bank2[1303], bank1[1303], bank0[1303]} = 32'h0;
    {bank3[1304], bank2[1304], bank1[1304], bank0[1304]} = 32'h0;
    {bank3[1305], bank2[1305], bank1[1305], bank0[1305]} = 32'h0;
    {bank3[1306], bank2[1306], bank1[1306], bank0[1306]} = 32'h0;
    {bank3[1307], bank2[1307], bank1[1307], bank0[1307]} = 32'h0;
    {bank3[1308], bank2[1308], bank1[1308], bank0[1308]} = 32'h0;
    {bank3[1309], bank2[1309], bank1[1309], bank0[1309]} = 32'h0;
    {bank3[1310], bank2[1310], bank1[1310], bank0[1310]} = 32'h0;
    {bank3[1311], bank2[1311], bank1[1311], bank0[1311]} = 32'h0;
    {bank3[1312], bank2[1312], bank1[1312], bank0[1312]} = 32'h0;
    {bank3[1313], bank2[1313], bank1[1313], bank0[1313]} = 32'h0;
    {bank3[1314], bank2[1314], bank1[1314], bank0[1314]} = 32'h0;
    {bank3[1315], bank2[1315], bank1[1315], bank0[1315]} = 32'h0;
    {bank3[1316], bank2[1316], bank1[1316], bank0[1316]} = 32'h0;
    {bank3[1317], bank2[1317], bank1[1317], bank0[1317]} = 32'h0;
    {bank3[1318], bank2[1318], bank1[1318], bank0[1318]} = 32'h0;
    {bank3[1319], bank2[1319], bank1[1319], bank0[1319]} = 32'h0;
    {bank3[1320], bank2[1320], bank1[1320], bank0[1320]} = 32'h0;
    {bank3[1321], bank2[1321], bank1[1321], bank0[1321]} = 32'h0;
    {bank3[1322], bank2[1322], bank1[1322], bank0[1322]} = 32'h0;
    {bank3[1323], bank2[1323], bank1[1323], bank0[1323]} = 32'h0;
    {bank3[1324], bank2[1324], bank1[1324], bank0[1324]} = 32'h0;
    {bank3[1325], bank2[1325], bank1[1325], bank0[1325]} = 32'h0;
    {bank3[1326], bank2[1326], bank1[1326], bank0[1326]} = 32'h0;
    {bank3[1327], bank2[1327], bank1[1327], bank0[1327]} = 32'h0;
    {bank3[1328], bank2[1328], bank1[1328], bank0[1328]} = 32'h0;
    {bank3[1329], bank2[1329], bank1[1329], bank0[1329]} = 32'h0;
    {bank3[1330], bank2[1330], bank1[1330], bank0[1330]} = 32'h0;
    {bank3[1331], bank2[1331], bank1[1331], bank0[1331]} = 32'h0;
    {bank3[1332], bank2[1332], bank1[1332], bank0[1332]} = 32'h0;
    {bank3[1333], bank2[1333], bank1[1333], bank0[1333]} = 32'h0;
    {bank3[1334], bank2[1334], bank1[1334], bank0[1334]} = 32'h0;
    {bank3[1335], bank2[1335], bank1[1335], bank0[1335]} = 32'h0;
    {bank3[1336], bank2[1336], bank1[1336], bank0[1336]} = 32'h0;
    {bank3[1337], bank2[1337], bank1[1337], bank0[1337]} = 32'h0;
    {bank3[1338], bank2[1338], bank1[1338], bank0[1338]} = 32'h0;
    {bank3[1339], bank2[1339], bank1[1339], bank0[1339]} = 32'h0;
    {bank3[1340], bank2[1340], bank1[1340], bank0[1340]} = 32'h0;
    {bank3[1341], bank2[1341], bank1[1341], bank0[1341]} = 32'h0;
    {bank3[1342], bank2[1342], bank1[1342], bank0[1342]} = 32'h0;
    {bank3[1343], bank2[1343], bank1[1343], bank0[1343]} = 32'h0;
    {bank3[1344], bank2[1344], bank1[1344], bank0[1344]} = 32'h0;
    {bank3[1345], bank2[1345], bank1[1345], bank0[1345]} = 32'h0;
    {bank3[1346], bank2[1346], bank1[1346], bank0[1346]} = 32'h0;
    {bank3[1347], bank2[1347], bank1[1347], bank0[1347]} = 32'h0;
    {bank3[1348], bank2[1348], bank1[1348], bank0[1348]} = 32'h0;
    {bank3[1349], bank2[1349], bank1[1349], bank0[1349]} = 32'h0;
    {bank3[1350], bank2[1350], bank1[1350], bank0[1350]} = 32'h0;
    {bank3[1351], bank2[1351], bank1[1351], bank0[1351]} = 32'h0;
    {bank3[1352], bank2[1352], bank1[1352], bank0[1352]} = 32'h0;
    {bank3[1353], bank2[1353], bank1[1353], bank0[1353]} = 32'h0;
    {bank3[1354], bank2[1354], bank1[1354], bank0[1354]} = 32'h0;
    {bank3[1355], bank2[1355], bank1[1355], bank0[1355]} = 32'h0;
    {bank3[1356], bank2[1356], bank1[1356], bank0[1356]} = 32'h0;
    {bank3[1357], bank2[1357], bank1[1357], bank0[1357]} = 32'h0;
    {bank3[1358], bank2[1358], bank1[1358], bank0[1358]} = 32'h0;
    {bank3[1359], bank2[1359], bank1[1359], bank0[1359]} = 32'h0;
    {bank3[1360], bank2[1360], bank1[1360], bank0[1360]} = 32'h0;
    {bank3[1361], bank2[1361], bank1[1361], bank0[1361]} = 32'h0;
    {bank3[1362], bank2[1362], bank1[1362], bank0[1362]} = 32'h0;
    {bank3[1363], bank2[1363], bank1[1363], bank0[1363]} = 32'h0;
    {bank3[1364], bank2[1364], bank1[1364], bank0[1364]} = 32'h0;
    {bank3[1365], bank2[1365], bank1[1365], bank0[1365]} = 32'h0;
    {bank3[1366], bank2[1366], bank1[1366], bank0[1366]} = 32'h0;
    {bank3[1367], bank2[1367], bank1[1367], bank0[1367]} = 32'h0;
    {bank3[1368], bank2[1368], bank1[1368], bank0[1368]} = 32'h0;
    {bank3[1369], bank2[1369], bank1[1369], bank0[1369]} = 32'h0;
    {bank3[1370], bank2[1370], bank1[1370], bank0[1370]} = 32'h0;
    {bank3[1371], bank2[1371], bank1[1371], bank0[1371]} = 32'h0;
    {bank3[1372], bank2[1372], bank1[1372], bank0[1372]} = 32'h0;
    {bank3[1373], bank2[1373], bank1[1373], bank0[1373]} = 32'h0;
    {bank3[1374], bank2[1374], bank1[1374], bank0[1374]} = 32'h0;
    {bank3[1375], bank2[1375], bank1[1375], bank0[1375]} = 32'h0;
    {bank3[1376], bank2[1376], bank1[1376], bank0[1376]} = 32'h0;
    {bank3[1377], bank2[1377], bank1[1377], bank0[1377]} = 32'h0;
    {bank3[1378], bank2[1378], bank1[1378], bank0[1378]} = 32'h0;
    {bank3[1379], bank2[1379], bank1[1379], bank0[1379]} = 32'h0;
    {bank3[1380], bank2[1380], bank1[1380], bank0[1380]} = 32'h0;
    {bank3[1381], bank2[1381], bank1[1381], bank0[1381]} = 32'h0;
    {bank3[1382], bank2[1382], bank1[1382], bank0[1382]} = 32'h0;
    {bank3[1383], bank2[1383], bank1[1383], bank0[1383]} = 32'h0;
    {bank3[1384], bank2[1384], bank1[1384], bank0[1384]} = 32'h0;
    {bank3[1385], bank2[1385], bank1[1385], bank0[1385]} = 32'h0;
    {bank3[1386], bank2[1386], bank1[1386], bank0[1386]} = 32'h0;
    {bank3[1387], bank2[1387], bank1[1387], bank0[1387]} = 32'h0;
    {bank3[1388], bank2[1388], bank1[1388], bank0[1388]} = 32'h0;
    {bank3[1389], bank2[1389], bank1[1389], bank0[1389]} = 32'h0;
    {bank3[1390], bank2[1390], bank1[1390], bank0[1390]} = 32'h0;
    {bank3[1391], bank2[1391], bank1[1391], bank0[1391]} = 32'h0;
    {bank3[1392], bank2[1392], bank1[1392], bank0[1392]} = 32'h0;
    {bank3[1393], bank2[1393], bank1[1393], bank0[1393]} = 32'h0;
    {bank3[1394], bank2[1394], bank1[1394], bank0[1394]} = 32'h0;
    {bank3[1395], bank2[1395], bank1[1395], bank0[1395]} = 32'h0;
    {bank3[1396], bank2[1396], bank1[1396], bank0[1396]} = 32'h0;
    {bank3[1397], bank2[1397], bank1[1397], bank0[1397]} = 32'h0;
    {bank3[1398], bank2[1398], bank1[1398], bank0[1398]} = 32'h0;
    {bank3[1399], bank2[1399], bank1[1399], bank0[1399]} = 32'h0;
    {bank3[1400], bank2[1400], bank1[1400], bank0[1400]} = 32'h0;
    {bank3[1401], bank2[1401], bank1[1401], bank0[1401]} = 32'h0;
    {bank3[1402], bank2[1402], bank1[1402], bank0[1402]} = 32'h0;
    {bank3[1403], bank2[1403], bank1[1403], bank0[1403]} = 32'h0;
    {bank3[1404], bank2[1404], bank1[1404], bank0[1404]} = 32'h0;
    {bank3[1405], bank2[1405], bank1[1405], bank0[1405]} = 32'h0;
    {bank3[1406], bank2[1406], bank1[1406], bank0[1406]} = 32'h0;
    {bank3[1407], bank2[1407], bank1[1407], bank0[1407]} = 32'h0;
    {bank3[1408], bank2[1408], bank1[1408], bank0[1408]} = 32'h0;
    {bank3[1409], bank2[1409], bank1[1409], bank0[1409]} = 32'h0;
    {bank3[1410], bank2[1410], bank1[1410], bank0[1410]} = 32'h0;
    {bank3[1411], bank2[1411], bank1[1411], bank0[1411]} = 32'h0;
    {bank3[1412], bank2[1412], bank1[1412], bank0[1412]} = 32'h0;
    {bank3[1413], bank2[1413], bank1[1413], bank0[1413]} = 32'h0;
    {bank3[1414], bank2[1414], bank1[1414], bank0[1414]} = 32'h0;
    {bank3[1415], bank2[1415], bank1[1415], bank0[1415]} = 32'h0;
    {bank3[1416], bank2[1416], bank1[1416], bank0[1416]} = 32'h0;
    {bank3[1417], bank2[1417], bank1[1417], bank0[1417]} = 32'h0;
    {bank3[1418], bank2[1418], bank1[1418], bank0[1418]} = 32'h0;
    {bank3[1419], bank2[1419], bank1[1419], bank0[1419]} = 32'h0;
    {bank3[1420], bank2[1420], bank1[1420], bank0[1420]} = 32'h0;
    {bank3[1421], bank2[1421], bank1[1421], bank0[1421]} = 32'h0;
    {bank3[1422], bank2[1422], bank1[1422], bank0[1422]} = 32'h0;
    {bank3[1423], bank2[1423], bank1[1423], bank0[1423]} = 32'h0;
    {bank3[1424], bank2[1424], bank1[1424], bank0[1424]} = 32'h0;
    {bank3[1425], bank2[1425], bank1[1425], bank0[1425]} = 32'h0;
    {bank3[1426], bank2[1426], bank1[1426], bank0[1426]} = 32'h0;
    {bank3[1427], bank2[1427], bank1[1427], bank0[1427]} = 32'h0;
    {bank3[1428], bank2[1428], bank1[1428], bank0[1428]} = 32'h0;
    {bank3[1429], bank2[1429], bank1[1429], bank0[1429]} = 32'h0;
    {bank3[1430], bank2[1430], bank1[1430], bank0[1430]} = 32'h0;
    {bank3[1431], bank2[1431], bank1[1431], bank0[1431]} = 32'h0;
    {bank3[1432], bank2[1432], bank1[1432], bank0[1432]} = 32'h0;
    {bank3[1433], bank2[1433], bank1[1433], bank0[1433]} = 32'h0;
    {bank3[1434], bank2[1434], bank1[1434], bank0[1434]} = 32'h0;
    {bank3[1435], bank2[1435], bank1[1435], bank0[1435]} = 32'h0;
    {bank3[1436], bank2[1436], bank1[1436], bank0[1436]} = 32'h0;
    {bank3[1437], bank2[1437], bank1[1437], bank0[1437]} = 32'h0;
    {bank3[1438], bank2[1438], bank1[1438], bank0[1438]} = 32'h0;
    {bank3[1439], bank2[1439], bank1[1439], bank0[1439]} = 32'h0;
    {bank3[1440], bank2[1440], bank1[1440], bank0[1440]} = 32'h0;
    {bank3[1441], bank2[1441], bank1[1441], bank0[1441]} = 32'h0;
    {bank3[1442], bank2[1442], bank1[1442], bank0[1442]} = 32'h0;
    {bank3[1443], bank2[1443], bank1[1443], bank0[1443]} = 32'h0;
    {bank3[1444], bank2[1444], bank1[1444], bank0[1444]} = 32'h0;
    {bank3[1445], bank2[1445], bank1[1445], bank0[1445]} = 32'h0;
    {bank3[1446], bank2[1446], bank1[1446], bank0[1446]} = 32'h0;
    {bank3[1447], bank2[1447], bank1[1447], bank0[1447]} = 32'h0;
    {bank3[1448], bank2[1448], bank1[1448], bank0[1448]} = 32'h0;
    {bank3[1449], bank2[1449], bank1[1449], bank0[1449]} = 32'h0;
    {bank3[1450], bank2[1450], bank1[1450], bank0[1450]} = 32'h0;
    {bank3[1451], bank2[1451], bank1[1451], bank0[1451]} = 32'h0;
    {bank3[1452], bank2[1452], bank1[1452], bank0[1452]} = 32'h0;
    {bank3[1453], bank2[1453], bank1[1453], bank0[1453]} = 32'h0;
    {bank3[1454], bank2[1454], bank1[1454], bank0[1454]} = 32'h0;
    {bank3[1455], bank2[1455], bank1[1455], bank0[1455]} = 32'h0;
    {bank3[1456], bank2[1456], bank1[1456], bank0[1456]} = 32'h0;
    {bank3[1457], bank2[1457], bank1[1457], bank0[1457]} = 32'h0;
    {bank3[1458], bank2[1458], bank1[1458], bank0[1458]} = 32'h0;
    {bank3[1459], bank2[1459], bank1[1459], bank0[1459]} = 32'h0;
    {bank3[1460], bank2[1460], bank1[1460], bank0[1460]} = 32'h0;
    {bank3[1461], bank2[1461], bank1[1461], bank0[1461]} = 32'h0;
    {bank3[1462], bank2[1462], bank1[1462], bank0[1462]} = 32'h0;
    {bank3[1463], bank2[1463], bank1[1463], bank0[1463]} = 32'h0;
    {bank3[1464], bank2[1464], bank1[1464], bank0[1464]} = 32'h0;
    {bank3[1465], bank2[1465], bank1[1465], bank0[1465]} = 32'h0;
    {bank3[1466], bank2[1466], bank1[1466], bank0[1466]} = 32'h0;
    {bank3[1467], bank2[1467], bank1[1467], bank0[1467]} = 32'h0;
    {bank3[1468], bank2[1468], bank1[1468], bank0[1468]} = 32'h0;
    {bank3[1469], bank2[1469], bank1[1469], bank0[1469]} = 32'h0;
    {bank3[1470], bank2[1470], bank1[1470], bank0[1470]} = 32'h0;
    {bank3[1471], bank2[1471], bank1[1471], bank0[1471]} = 32'h0;
    {bank3[1472], bank2[1472], bank1[1472], bank0[1472]} = 32'h0;
    {bank3[1473], bank2[1473], bank1[1473], bank0[1473]} = 32'h0;
    {bank3[1474], bank2[1474], bank1[1474], bank0[1474]} = 32'h0;
    {bank3[1475], bank2[1475], bank1[1475], bank0[1475]} = 32'h0;
    {bank3[1476], bank2[1476], bank1[1476], bank0[1476]} = 32'h0;
    {bank3[1477], bank2[1477], bank1[1477], bank0[1477]} = 32'h0;
    {bank3[1478], bank2[1478], bank1[1478], bank0[1478]} = 32'h0;
    {bank3[1479], bank2[1479], bank1[1479], bank0[1479]} = 32'h0;
    {bank3[1480], bank2[1480], bank1[1480], bank0[1480]} = 32'h0;
    {bank3[1481], bank2[1481], bank1[1481], bank0[1481]} = 32'h0;
    {bank3[1482], bank2[1482], bank1[1482], bank0[1482]} = 32'h0;
    {bank3[1483], bank2[1483], bank1[1483], bank0[1483]} = 32'h0;
    {bank3[1484], bank2[1484], bank1[1484], bank0[1484]} = 32'h0;
    {bank3[1485], bank2[1485], bank1[1485], bank0[1485]} = 32'h0;
    {bank3[1486], bank2[1486], bank1[1486], bank0[1486]} = 32'h0;
    {bank3[1487], bank2[1487], bank1[1487], bank0[1487]} = 32'h0;
    {bank3[1488], bank2[1488], bank1[1488], bank0[1488]} = 32'h0;
    {bank3[1489], bank2[1489], bank1[1489], bank0[1489]} = 32'h0;
    {bank3[1490], bank2[1490], bank1[1490], bank0[1490]} = 32'h0;
    {bank3[1491], bank2[1491], bank1[1491], bank0[1491]} = 32'h0;
    {bank3[1492], bank2[1492], bank1[1492], bank0[1492]} = 32'h0;
    {bank3[1493], bank2[1493], bank1[1493], bank0[1493]} = 32'h0;
    {bank3[1494], bank2[1494], bank1[1494], bank0[1494]} = 32'h0;
    {bank3[1495], bank2[1495], bank1[1495], bank0[1495]} = 32'h0;
    {bank3[1496], bank2[1496], bank1[1496], bank0[1496]} = 32'h0;
    {bank3[1497], bank2[1497], bank1[1497], bank0[1497]} = 32'h0;
    {bank3[1498], bank2[1498], bank1[1498], bank0[1498]} = 32'h0;
    {bank3[1499], bank2[1499], bank1[1499], bank0[1499]} = 32'h0;
    {bank3[1500], bank2[1500], bank1[1500], bank0[1500]} = 32'h0;
    {bank3[1501], bank2[1501], bank1[1501], bank0[1501]} = 32'h0;
    {bank3[1502], bank2[1502], bank1[1502], bank0[1502]} = 32'h0;
    {bank3[1503], bank2[1503], bank1[1503], bank0[1503]} = 32'h0;
    {bank3[1504], bank2[1504], bank1[1504], bank0[1504]} = 32'h0;
    {bank3[1505], bank2[1505], bank1[1505], bank0[1505]} = 32'h0;
    {bank3[1506], bank2[1506], bank1[1506], bank0[1506]} = 32'h0;
    {bank3[1507], bank2[1507], bank1[1507], bank0[1507]} = 32'h0;
    {bank3[1508], bank2[1508], bank1[1508], bank0[1508]} = 32'h0;
    {bank3[1509], bank2[1509], bank1[1509], bank0[1509]} = 32'h0;
    {bank3[1510], bank2[1510], bank1[1510], bank0[1510]} = 32'h0;
    {bank3[1511], bank2[1511], bank1[1511], bank0[1511]} = 32'h0;
    {bank3[1512], bank2[1512], bank1[1512], bank0[1512]} = 32'h0;
    {bank3[1513], bank2[1513], bank1[1513], bank0[1513]} = 32'h0;
    {bank3[1514], bank2[1514], bank1[1514], bank0[1514]} = 32'h0;
    {bank3[1515], bank2[1515], bank1[1515], bank0[1515]} = 32'h0;
    {bank3[1516], bank2[1516], bank1[1516], bank0[1516]} = 32'h0;
    {bank3[1517], bank2[1517], bank1[1517], bank0[1517]} = 32'h0;
    {bank3[1518], bank2[1518], bank1[1518], bank0[1518]} = 32'h0;
    {bank3[1519], bank2[1519], bank1[1519], bank0[1519]} = 32'h0;
    {bank3[1520], bank2[1520], bank1[1520], bank0[1520]} = 32'h0;
    {bank3[1521], bank2[1521], bank1[1521], bank0[1521]} = 32'h0;
    {bank3[1522], bank2[1522], bank1[1522], bank0[1522]} = 32'h0;
    {bank3[1523], bank2[1523], bank1[1523], bank0[1523]} = 32'h0;
    {bank3[1524], bank2[1524], bank1[1524], bank0[1524]} = 32'h0;
    {bank3[1525], bank2[1525], bank1[1525], bank0[1525]} = 32'h0;
    {bank3[1526], bank2[1526], bank1[1526], bank0[1526]} = 32'h0;
    {bank3[1527], bank2[1527], bank1[1527], bank0[1527]} = 32'h0;
    {bank3[1528], bank2[1528], bank1[1528], bank0[1528]} = 32'h0;
    {bank3[1529], bank2[1529], bank1[1529], bank0[1529]} = 32'h0;
    {bank3[1530], bank2[1530], bank1[1530], bank0[1530]} = 32'h0;
    {bank3[1531], bank2[1531], bank1[1531], bank0[1531]} = 32'h0;
    {bank3[1532], bank2[1532], bank1[1532], bank0[1532]} = 32'h0;
    {bank3[1533], bank2[1533], bank1[1533], bank0[1533]} = 32'h0;
    {bank3[1534], bank2[1534], bank1[1534], bank0[1534]} = 32'h0;
    {bank3[1535], bank2[1535], bank1[1535], bank0[1535]} = 32'h0;
    {bank3[1536], bank2[1536], bank1[1536], bank0[1536]} = 32'h0;
    {bank3[1537], bank2[1537], bank1[1537], bank0[1537]} = 32'h0;
    {bank3[1538], bank2[1538], bank1[1538], bank0[1538]} = 32'h0;
    {bank3[1539], bank2[1539], bank1[1539], bank0[1539]} = 32'h0;
    {bank3[1540], bank2[1540], bank1[1540], bank0[1540]} = 32'h0;
    {bank3[1541], bank2[1541], bank1[1541], bank0[1541]} = 32'h0;
    {bank3[1542], bank2[1542], bank1[1542], bank0[1542]} = 32'h0;
    {bank3[1543], bank2[1543], bank1[1543], bank0[1543]} = 32'h0;
    {bank3[1544], bank2[1544], bank1[1544], bank0[1544]} = 32'h0;
    {bank3[1545], bank2[1545], bank1[1545], bank0[1545]} = 32'h0;
    {bank3[1546], bank2[1546], bank1[1546], bank0[1546]} = 32'h0;
    {bank3[1547], bank2[1547], bank1[1547], bank0[1547]} = 32'h0;
    {bank3[1548], bank2[1548], bank1[1548], bank0[1548]} = 32'h0;
    {bank3[1549], bank2[1549], bank1[1549], bank0[1549]} = 32'h0;
    {bank3[1550], bank2[1550], bank1[1550], bank0[1550]} = 32'h0;
    {bank3[1551], bank2[1551], bank1[1551], bank0[1551]} = 32'h0;
    {bank3[1552], bank2[1552], bank1[1552], bank0[1552]} = 32'h0;
    {bank3[1553], bank2[1553], bank1[1553], bank0[1553]} = 32'h0;
    {bank3[1554], bank2[1554], bank1[1554], bank0[1554]} = 32'h0;
    {bank3[1555], bank2[1555], bank1[1555], bank0[1555]} = 32'h0;
    {bank3[1556], bank2[1556], bank1[1556], bank0[1556]} = 32'h0;
    {bank3[1557], bank2[1557], bank1[1557], bank0[1557]} = 32'h0;
    {bank3[1558], bank2[1558], bank1[1558], bank0[1558]} = 32'h0;
    {bank3[1559], bank2[1559], bank1[1559], bank0[1559]} = 32'h0;
    {bank3[1560], bank2[1560], bank1[1560], bank0[1560]} = 32'h0;
    {bank3[1561], bank2[1561], bank1[1561], bank0[1561]} = 32'h0;
    {bank3[1562], bank2[1562], bank1[1562], bank0[1562]} = 32'h0;
    {bank3[1563], bank2[1563], bank1[1563], bank0[1563]} = 32'h0;
    {bank3[1564], bank2[1564], bank1[1564], bank0[1564]} = 32'h0;
    {bank3[1565], bank2[1565], bank1[1565], bank0[1565]} = 32'h0;
    {bank3[1566], bank2[1566], bank1[1566], bank0[1566]} = 32'h0;
    {bank3[1567], bank2[1567], bank1[1567], bank0[1567]} = 32'h0;
    {bank3[1568], bank2[1568], bank1[1568], bank0[1568]} = 32'h0;
    {bank3[1569], bank2[1569], bank1[1569], bank0[1569]} = 32'h0;
    {bank3[1570], bank2[1570], bank1[1570], bank0[1570]} = 32'h0;
    {bank3[1571], bank2[1571], bank1[1571], bank0[1571]} = 32'h0;
    {bank3[1572], bank2[1572], bank1[1572], bank0[1572]} = 32'h0;
    {bank3[1573], bank2[1573], bank1[1573], bank0[1573]} = 32'h0;
    {bank3[1574], bank2[1574], bank1[1574], bank0[1574]} = 32'h0;
    {bank3[1575], bank2[1575], bank1[1575], bank0[1575]} = 32'h0;
    {bank3[1576], bank2[1576], bank1[1576], bank0[1576]} = 32'h0;
    {bank3[1577], bank2[1577], bank1[1577], bank0[1577]} = 32'h0;
    {bank3[1578], bank2[1578], bank1[1578], bank0[1578]} = 32'h0;
    {bank3[1579], bank2[1579], bank1[1579], bank0[1579]} = 32'h0;
    {bank3[1580], bank2[1580], bank1[1580], bank0[1580]} = 32'h0;
    {bank3[1581], bank2[1581], bank1[1581], bank0[1581]} = 32'h0;
    {bank3[1582], bank2[1582], bank1[1582], bank0[1582]} = 32'h0;
    {bank3[1583], bank2[1583], bank1[1583], bank0[1583]} = 32'h0;
    {bank3[1584], bank2[1584], bank1[1584], bank0[1584]} = 32'h0;
    {bank3[1585], bank2[1585], bank1[1585], bank0[1585]} = 32'h0;
    {bank3[1586], bank2[1586], bank1[1586], bank0[1586]} = 32'h0;
    {bank3[1587], bank2[1587], bank1[1587], bank0[1587]} = 32'h0;
    {bank3[1588], bank2[1588], bank1[1588], bank0[1588]} = 32'h0;
    {bank3[1589], bank2[1589], bank1[1589], bank0[1589]} = 32'h0;
    {bank3[1590], bank2[1590], bank1[1590], bank0[1590]} = 32'h0;
    {bank3[1591], bank2[1591], bank1[1591], bank0[1591]} = 32'h0;
    {bank3[1592], bank2[1592], bank1[1592], bank0[1592]} = 32'h0;
    {bank3[1593], bank2[1593], bank1[1593], bank0[1593]} = 32'h0;
    {bank3[1594], bank2[1594], bank1[1594], bank0[1594]} = 32'h0;
    {bank3[1595], bank2[1595], bank1[1595], bank0[1595]} = 32'h0;
    {bank3[1596], bank2[1596], bank1[1596], bank0[1596]} = 32'h0;
    {bank3[1597], bank2[1597], bank1[1597], bank0[1597]} = 32'h0;
    {bank3[1598], bank2[1598], bank1[1598], bank0[1598]} = 32'h0;
    {bank3[1599], bank2[1599], bank1[1599], bank0[1599]} = 32'h0;
    {bank3[1600], bank2[1600], bank1[1600], bank0[1600]} = 32'h0;
    {bank3[1601], bank2[1601], bank1[1601], bank0[1601]} = 32'h0;
    {bank3[1602], bank2[1602], bank1[1602], bank0[1602]} = 32'h0;
    {bank3[1603], bank2[1603], bank1[1603], bank0[1603]} = 32'h0;
    {bank3[1604], bank2[1604], bank1[1604], bank0[1604]} = 32'h0;
    {bank3[1605], bank2[1605], bank1[1605], bank0[1605]} = 32'h0;
    {bank3[1606], bank2[1606], bank1[1606], bank0[1606]} = 32'h0;
    {bank3[1607], bank2[1607], bank1[1607], bank0[1607]} = 32'h0;
    {bank3[1608], bank2[1608], bank1[1608], bank0[1608]} = 32'h0;
    {bank3[1609], bank2[1609], bank1[1609], bank0[1609]} = 32'h0;
    {bank3[1610], bank2[1610], bank1[1610], bank0[1610]} = 32'h0;
    {bank3[1611], bank2[1611], bank1[1611], bank0[1611]} = 32'h0;
    {bank3[1612], bank2[1612], bank1[1612], bank0[1612]} = 32'h0;
    {bank3[1613], bank2[1613], bank1[1613], bank0[1613]} = 32'h0;
    {bank3[1614], bank2[1614], bank1[1614], bank0[1614]} = 32'h0;
    {bank3[1615], bank2[1615], bank1[1615], bank0[1615]} = 32'h0;
    {bank3[1616], bank2[1616], bank1[1616], bank0[1616]} = 32'h0;
    {bank3[1617], bank2[1617], bank1[1617], bank0[1617]} = 32'h0;
    {bank3[1618], bank2[1618], bank1[1618], bank0[1618]} = 32'h0;
    {bank3[1619], bank2[1619], bank1[1619], bank0[1619]} = 32'h0;
    {bank3[1620], bank2[1620], bank1[1620], bank0[1620]} = 32'h0;
    {bank3[1621], bank2[1621], bank1[1621], bank0[1621]} = 32'h0;
    {bank3[1622], bank2[1622], bank1[1622], bank0[1622]} = 32'h0;
    {bank3[1623], bank2[1623], bank1[1623], bank0[1623]} = 32'h0;
    {bank3[1624], bank2[1624], bank1[1624], bank0[1624]} = 32'h0;
    {bank3[1625], bank2[1625], bank1[1625], bank0[1625]} = 32'h0;
    {bank3[1626], bank2[1626], bank1[1626], bank0[1626]} = 32'h0;
    {bank3[1627], bank2[1627], bank1[1627], bank0[1627]} = 32'h0;
    {bank3[1628], bank2[1628], bank1[1628], bank0[1628]} = 32'h0;
    {bank3[1629], bank2[1629], bank1[1629], bank0[1629]} = 32'h0;
    {bank3[1630], bank2[1630], bank1[1630], bank0[1630]} = 32'h0;
    {bank3[1631], bank2[1631], bank1[1631], bank0[1631]} = 32'h0;
    {bank3[1632], bank2[1632], bank1[1632], bank0[1632]} = 32'h0;
    {bank3[1633], bank2[1633], bank1[1633], bank0[1633]} = 32'h0;
    {bank3[1634], bank2[1634], bank1[1634], bank0[1634]} = 32'h0;
    {bank3[1635], bank2[1635], bank1[1635], bank0[1635]} = 32'h0;
    {bank3[1636], bank2[1636], bank1[1636], bank0[1636]} = 32'h0;
    {bank3[1637], bank2[1637], bank1[1637], bank0[1637]} = 32'h0;
    {bank3[1638], bank2[1638], bank1[1638], bank0[1638]} = 32'h0;
    {bank3[1639], bank2[1639], bank1[1639], bank0[1639]} = 32'h0;
    {bank3[1640], bank2[1640], bank1[1640], bank0[1640]} = 32'h0;
    {bank3[1641], bank2[1641], bank1[1641], bank0[1641]} = 32'h0;
    {bank3[1642], bank2[1642], bank1[1642], bank0[1642]} = 32'h0;
    {bank3[1643], bank2[1643], bank1[1643], bank0[1643]} = 32'h0;
    {bank3[1644], bank2[1644], bank1[1644], bank0[1644]} = 32'h0;
    {bank3[1645], bank2[1645], bank1[1645], bank0[1645]} = 32'h0;
    {bank3[1646], bank2[1646], bank1[1646], bank0[1646]} = 32'h0;
    {bank3[1647], bank2[1647], bank1[1647], bank0[1647]} = 32'h0;
    {bank3[1648], bank2[1648], bank1[1648], bank0[1648]} = 32'h0;
    {bank3[1649], bank2[1649], bank1[1649], bank0[1649]} = 32'h0;
    {bank3[1650], bank2[1650], bank1[1650], bank0[1650]} = 32'h0;
    {bank3[1651], bank2[1651], bank1[1651], bank0[1651]} = 32'h0;
    {bank3[1652], bank2[1652], bank1[1652], bank0[1652]} = 32'h0;
    {bank3[1653], bank2[1653], bank1[1653], bank0[1653]} = 32'h0;
    {bank3[1654], bank2[1654], bank1[1654], bank0[1654]} = 32'h0;
    {bank3[1655], bank2[1655], bank1[1655], bank0[1655]} = 32'h0;
    {bank3[1656], bank2[1656], bank1[1656], bank0[1656]} = 32'h0;
    {bank3[1657], bank2[1657], bank1[1657], bank0[1657]} = 32'h0;
    {bank3[1658], bank2[1658], bank1[1658], bank0[1658]} = 32'h0;
    {bank3[1659], bank2[1659], bank1[1659], bank0[1659]} = 32'h0;
    {bank3[1660], bank2[1660], bank1[1660], bank0[1660]} = 32'h0;
    {bank3[1661], bank2[1661], bank1[1661], bank0[1661]} = 32'h0;
    {bank3[1662], bank2[1662], bank1[1662], bank0[1662]} = 32'h0;
    {bank3[1663], bank2[1663], bank1[1663], bank0[1663]} = 32'h0;
    {bank3[1664], bank2[1664], bank1[1664], bank0[1664]} = 32'h0;
    {bank3[1665], bank2[1665], bank1[1665], bank0[1665]} = 32'h0;
    {bank3[1666], bank2[1666], bank1[1666], bank0[1666]} = 32'h0;
    {bank3[1667], bank2[1667], bank1[1667], bank0[1667]} = 32'h0;
    {bank3[1668], bank2[1668], bank1[1668], bank0[1668]} = 32'h0;
    {bank3[1669], bank2[1669], bank1[1669], bank0[1669]} = 32'h0;
    {bank3[1670], bank2[1670], bank1[1670], bank0[1670]} = 32'h0;
    {bank3[1671], bank2[1671], bank1[1671], bank0[1671]} = 32'h0;
    {bank3[1672], bank2[1672], bank1[1672], bank0[1672]} = 32'h0;
    {bank3[1673], bank2[1673], bank1[1673], bank0[1673]} = 32'h0;
    {bank3[1674], bank2[1674], bank1[1674], bank0[1674]} = 32'h0;
    {bank3[1675], bank2[1675], bank1[1675], bank0[1675]} = 32'h0;
    {bank3[1676], bank2[1676], bank1[1676], bank0[1676]} = 32'h0;
    {bank3[1677], bank2[1677], bank1[1677], bank0[1677]} = 32'h0;
    {bank3[1678], bank2[1678], bank1[1678], bank0[1678]} = 32'h0;
    {bank3[1679], bank2[1679], bank1[1679], bank0[1679]} = 32'h0;
    {bank3[1680], bank2[1680], bank1[1680], bank0[1680]} = 32'h0;
    {bank3[1681], bank2[1681], bank1[1681], bank0[1681]} = 32'h0;
    {bank3[1682], bank2[1682], bank1[1682], bank0[1682]} = 32'h0;
    {bank3[1683], bank2[1683], bank1[1683], bank0[1683]} = 32'h0;
    {bank3[1684], bank2[1684], bank1[1684], bank0[1684]} = 32'h0;
    {bank3[1685], bank2[1685], bank1[1685], bank0[1685]} = 32'h0;
    {bank3[1686], bank2[1686], bank1[1686], bank0[1686]} = 32'h0;
    {bank3[1687], bank2[1687], bank1[1687], bank0[1687]} = 32'h0;
    {bank3[1688], bank2[1688], bank1[1688], bank0[1688]} = 32'h0;
    {bank3[1689], bank2[1689], bank1[1689], bank0[1689]} = 32'h0;
    {bank3[1690], bank2[1690], bank1[1690], bank0[1690]} = 32'h0;
    {bank3[1691], bank2[1691], bank1[1691], bank0[1691]} = 32'h0;
    {bank3[1692], bank2[1692], bank1[1692], bank0[1692]} = 32'h0;
    {bank3[1693], bank2[1693], bank1[1693], bank0[1693]} = 32'h0;
    {bank3[1694], bank2[1694], bank1[1694], bank0[1694]} = 32'h0;
    {bank3[1695], bank2[1695], bank1[1695], bank0[1695]} = 32'h0;
    {bank3[1696], bank2[1696], bank1[1696], bank0[1696]} = 32'h0;
    {bank3[1697], bank2[1697], bank1[1697], bank0[1697]} = 32'h0;
    {bank3[1698], bank2[1698], bank1[1698], bank0[1698]} = 32'h0;
    {bank3[1699], bank2[1699], bank1[1699], bank0[1699]} = 32'h0;
    {bank3[1700], bank2[1700], bank1[1700], bank0[1700]} = 32'h0;
    {bank3[1701], bank2[1701], bank1[1701], bank0[1701]} = 32'h0;
    {bank3[1702], bank2[1702], bank1[1702], bank0[1702]} = 32'h0;
    {bank3[1703], bank2[1703], bank1[1703], bank0[1703]} = 32'h0;
    {bank3[1704], bank2[1704], bank1[1704], bank0[1704]} = 32'h0;
    {bank3[1705], bank2[1705], bank1[1705], bank0[1705]} = 32'h0;
    {bank3[1706], bank2[1706], bank1[1706], bank0[1706]} = 32'h0;
    {bank3[1707], bank2[1707], bank1[1707], bank0[1707]} = 32'h0;
    {bank3[1708], bank2[1708], bank1[1708], bank0[1708]} = 32'h0;
    {bank3[1709], bank2[1709], bank1[1709], bank0[1709]} = 32'h0;
    {bank3[1710], bank2[1710], bank1[1710], bank0[1710]} = 32'h0;
    {bank3[1711], bank2[1711], bank1[1711], bank0[1711]} = 32'h0;
    {bank3[1712], bank2[1712], bank1[1712], bank0[1712]} = 32'h0;
    {bank3[1713], bank2[1713], bank1[1713], bank0[1713]} = 32'h0;
    {bank3[1714], bank2[1714], bank1[1714], bank0[1714]} = 32'h0;
    {bank3[1715], bank2[1715], bank1[1715], bank0[1715]} = 32'h0;
    {bank3[1716], bank2[1716], bank1[1716], bank0[1716]} = 32'h0;
    {bank3[1717], bank2[1717], bank1[1717], bank0[1717]} = 32'h0;
    {bank3[1718], bank2[1718], bank1[1718], bank0[1718]} = 32'h0;
    {bank3[1719], bank2[1719], bank1[1719], bank0[1719]} = 32'h0;
    {bank3[1720], bank2[1720], bank1[1720], bank0[1720]} = 32'h0;
    {bank3[1721], bank2[1721], bank1[1721], bank0[1721]} = 32'h0;
    {bank3[1722], bank2[1722], bank1[1722], bank0[1722]} = 32'h0;
    {bank3[1723], bank2[1723], bank1[1723], bank0[1723]} = 32'h0;
    {bank3[1724], bank2[1724], bank1[1724], bank0[1724]} = 32'h0;
    {bank3[1725], bank2[1725], bank1[1725], bank0[1725]} = 32'h0;
    {bank3[1726], bank2[1726], bank1[1726], bank0[1726]} = 32'h0;
    {bank3[1727], bank2[1727], bank1[1727], bank0[1727]} = 32'h0;
    {bank3[1728], bank2[1728], bank1[1728], bank0[1728]} = 32'h0;
    {bank3[1729], bank2[1729], bank1[1729], bank0[1729]} = 32'h0;
    {bank3[1730], bank2[1730], bank1[1730], bank0[1730]} = 32'h0;
    {bank3[1731], bank2[1731], bank1[1731], bank0[1731]} = 32'h0;
    {bank3[1732], bank2[1732], bank1[1732], bank0[1732]} = 32'h0;
    {bank3[1733], bank2[1733], bank1[1733], bank0[1733]} = 32'h0;
    {bank3[1734], bank2[1734], bank1[1734], bank0[1734]} = 32'h0;
    {bank3[1735], bank2[1735], bank1[1735], bank0[1735]} = 32'h0;
    {bank3[1736], bank2[1736], bank1[1736], bank0[1736]} = 32'h0;
    {bank3[1737], bank2[1737], bank1[1737], bank0[1737]} = 32'h0;
    {bank3[1738], bank2[1738], bank1[1738], bank0[1738]} = 32'h0;
    {bank3[1739], bank2[1739], bank1[1739], bank0[1739]} = 32'h0;
    {bank3[1740], bank2[1740], bank1[1740], bank0[1740]} = 32'h0;
    {bank3[1741], bank2[1741], bank1[1741], bank0[1741]} = 32'h0;
    {bank3[1742], bank2[1742], bank1[1742], bank0[1742]} = 32'h0;
    {bank3[1743], bank2[1743], bank1[1743], bank0[1743]} = 32'h0;
    {bank3[1744], bank2[1744], bank1[1744], bank0[1744]} = 32'h0;
    {bank3[1745], bank2[1745], bank1[1745], bank0[1745]} = 32'h0;
    {bank3[1746], bank2[1746], bank1[1746], bank0[1746]} = 32'h0;
    {bank3[1747], bank2[1747], bank1[1747], bank0[1747]} = 32'h0;
    {bank3[1748], bank2[1748], bank1[1748], bank0[1748]} = 32'h0;
    {bank3[1749], bank2[1749], bank1[1749], bank0[1749]} = 32'h0;
    {bank3[1750], bank2[1750], bank1[1750], bank0[1750]} = 32'h0;
    {bank3[1751], bank2[1751], bank1[1751], bank0[1751]} = 32'h0;
    {bank3[1752], bank2[1752], bank1[1752], bank0[1752]} = 32'h0;
    {bank3[1753], bank2[1753], bank1[1753], bank0[1753]} = 32'h0;
    {bank3[1754], bank2[1754], bank1[1754], bank0[1754]} = 32'h0;
    {bank3[1755], bank2[1755], bank1[1755], bank0[1755]} = 32'h0;
    {bank3[1756], bank2[1756], bank1[1756], bank0[1756]} = 32'h0;
    {bank3[1757], bank2[1757], bank1[1757], bank0[1757]} = 32'h0;
    {bank3[1758], bank2[1758], bank1[1758], bank0[1758]} = 32'h0;
    {bank3[1759], bank2[1759], bank1[1759], bank0[1759]} = 32'h0;
    {bank3[1760], bank2[1760], bank1[1760], bank0[1760]} = 32'h0;
    {bank3[1761], bank2[1761], bank1[1761], bank0[1761]} = 32'h0;
    {bank3[1762], bank2[1762], bank1[1762], bank0[1762]} = 32'h0;
    {bank3[1763], bank2[1763], bank1[1763], bank0[1763]} = 32'h0;
    {bank3[1764], bank2[1764], bank1[1764], bank0[1764]} = 32'h0;
    {bank3[1765], bank2[1765], bank1[1765], bank0[1765]} = 32'h0;
    {bank3[1766], bank2[1766], bank1[1766], bank0[1766]} = 32'h0;
    {bank3[1767], bank2[1767], bank1[1767], bank0[1767]} = 32'h0;
    {bank3[1768], bank2[1768], bank1[1768], bank0[1768]} = 32'h0;
    {bank3[1769], bank2[1769], bank1[1769], bank0[1769]} = 32'h0;
    {bank3[1770], bank2[1770], bank1[1770], bank0[1770]} = 32'h0;
    {bank3[1771], bank2[1771], bank1[1771], bank0[1771]} = 32'h0;
    {bank3[1772], bank2[1772], bank1[1772], bank0[1772]} = 32'h0;
    {bank3[1773], bank2[1773], bank1[1773], bank0[1773]} = 32'h0;
    {bank3[1774], bank2[1774], bank1[1774], bank0[1774]} = 32'h0;
    {bank3[1775], bank2[1775], bank1[1775], bank0[1775]} = 32'h0;
    {bank3[1776], bank2[1776], bank1[1776], bank0[1776]} = 32'h0;
    {bank3[1777], bank2[1777], bank1[1777], bank0[1777]} = 32'h0;
    {bank3[1778], bank2[1778], bank1[1778], bank0[1778]} = 32'h0;
    {bank3[1779], bank2[1779], bank1[1779], bank0[1779]} = 32'h0;
    {bank3[1780], bank2[1780], bank1[1780], bank0[1780]} = 32'h0;
    {bank3[1781], bank2[1781], bank1[1781], bank0[1781]} = 32'h0;
    {bank3[1782], bank2[1782], bank1[1782], bank0[1782]} = 32'h0;
    {bank3[1783], bank2[1783], bank1[1783], bank0[1783]} = 32'h0;
    {bank3[1784], bank2[1784], bank1[1784], bank0[1784]} = 32'h0;
    {bank3[1785], bank2[1785], bank1[1785], bank0[1785]} = 32'h0;
    {bank3[1786], bank2[1786], bank1[1786], bank0[1786]} = 32'h0;
    {bank3[1787], bank2[1787], bank1[1787], bank0[1787]} = 32'h0;
    {bank3[1788], bank2[1788], bank1[1788], bank0[1788]} = 32'h0;
    {bank3[1789], bank2[1789], bank1[1789], bank0[1789]} = 32'h0;
    {bank3[1790], bank2[1790], bank1[1790], bank0[1790]} = 32'h0;
    {bank3[1791], bank2[1791], bank1[1791], bank0[1791]} = 32'h0;
    {bank3[1792], bank2[1792], bank1[1792], bank0[1792]} = 32'h0;
    {bank3[1793], bank2[1793], bank1[1793], bank0[1793]} = 32'h0;
    {bank3[1794], bank2[1794], bank1[1794], bank0[1794]} = 32'h0;
    {bank3[1795], bank2[1795], bank1[1795], bank0[1795]} = 32'h0;
    {bank3[1796], bank2[1796], bank1[1796], bank0[1796]} = 32'h0;
    {bank3[1797], bank2[1797], bank1[1797], bank0[1797]} = 32'h0;
    {bank3[1798], bank2[1798], bank1[1798], bank0[1798]} = 32'h0;
    {bank3[1799], bank2[1799], bank1[1799], bank0[1799]} = 32'h0;
    {bank3[1800], bank2[1800], bank1[1800], bank0[1800]} = 32'h0;
    {bank3[1801], bank2[1801], bank1[1801], bank0[1801]} = 32'h0;
    {bank3[1802], bank2[1802], bank1[1802], bank0[1802]} = 32'h0;
    {bank3[1803], bank2[1803], bank1[1803], bank0[1803]} = 32'h0;
    {bank3[1804], bank2[1804], bank1[1804], bank0[1804]} = 32'h0;
    {bank3[1805], bank2[1805], bank1[1805], bank0[1805]} = 32'h0;
    {bank3[1806], bank2[1806], bank1[1806], bank0[1806]} = 32'h0;
    {bank3[1807], bank2[1807], bank1[1807], bank0[1807]} = 32'h0;
    {bank3[1808], bank2[1808], bank1[1808], bank0[1808]} = 32'h0;
    {bank3[1809], bank2[1809], bank1[1809], bank0[1809]} = 32'h0;
    {bank3[1810], bank2[1810], bank1[1810], bank0[1810]} = 32'h0;
    {bank3[1811], bank2[1811], bank1[1811], bank0[1811]} = 32'h0;
    {bank3[1812], bank2[1812], bank1[1812], bank0[1812]} = 32'h0;
    {bank3[1813], bank2[1813], bank1[1813], bank0[1813]} = 32'h0;
    {bank3[1814], bank2[1814], bank1[1814], bank0[1814]} = 32'h0;
    {bank3[1815], bank2[1815], bank1[1815], bank0[1815]} = 32'h0;
    {bank3[1816], bank2[1816], bank1[1816], bank0[1816]} = 32'h0;
    {bank3[1817], bank2[1817], bank1[1817], bank0[1817]} = 32'h0;
    {bank3[1818], bank2[1818], bank1[1818], bank0[1818]} = 32'h0;
    {bank3[1819], bank2[1819], bank1[1819], bank0[1819]} = 32'h0;
    {bank3[1820], bank2[1820], bank1[1820], bank0[1820]} = 32'h0;
    {bank3[1821], bank2[1821], bank1[1821], bank0[1821]} = 32'h0;
    {bank3[1822], bank2[1822], bank1[1822], bank0[1822]} = 32'h0;
    {bank3[1823], bank2[1823], bank1[1823], bank0[1823]} = 32'h0;
    {bank3[1824], bank2[1824], bank1[1824], bank0[1824]} = 32'h0;
    {bank3[1825], bank2[1825], bank1[1825], bank0[1825]} = 32'h0;
    {bank3[1826], bank2[1826], bank1[1826], bank0[1826]} = 32'h0;
    {bank3[1827], bank2[1827], bank1[1827], bank0[1827]} = 32'h0;
    {bank3[1828], bank2[1828], bank1[1828], bank0[1828]} = 32'h0;
    {bank3[1829], bank2[1829], bank1[1829], bank0[1829]} = 32'h0;
    {bank3[1830], bank2[1830], bank1[1830], bank0[1830]} = 32'h0;
    {bank3[1831], bank2[1831], bank1[1831], bank0[1831]} = 32'h0;
    {bank3[1832], bank2[1832], bank1[1832], bank0[1832]} = 32'h0;
    {bank3[1833], bank2[1833], bank1[1833], bank0[1833]} = 32'h0;
    {bank3[1834], bank2[1834], bank1[1834], bank0[1834]} = 32'h0;
    {bank3[1835], bank2[1835], bank1[1835], bank0[1835]} = 32'h0;
    {bank3[1836], bank2[1836], bank1[1836], bank0[1836]} = 32'h0;
    {bank3[1837], bank2[1837], bank1[1837], bank0[1837]} = 32'h0;
    {bank3[1838], bank2[1838], bank1[1838], bank0[1838]} = 32'h0;
    {bank3[1839], bank2[1839], bank1[1839], bank0[1839]} = 32'h0;
    {bank3[1840], bank2[1840], bank1[1840], bank0[1840]} = 32'h0;
    {bank3[1841], bank2[1841], bank1[1841], bank0[1841]} = 32'h0;
    {bank3[1842], bank2[1842], bank1[1842], bank0[1842]} = 32'h0;
    {bank3[1843], bank2[1843], bank1[1843], bank0[1843]} = 32'h0;
    {bank3[1844], bank2[1844], bank1[1844], bank0[1844]} = 32'h0;
    {bank3[1845], bank2[1845], bank1[1845], bank0[1845]} = 32'h0;
    {bank3[1846], bank2[1846], bank1[1846], bank0[1846]} = 32'h0;
    {bank3[1847], bank2[1847], bank1[1847], bank0[1847]} = 32'h0;
    {bank3[1848], bank2[1848], bank1[1848], bank0[1848]} = 32'h0;
    {bank3[1849], bank2[1849], bank1[1849], bank0[1849]} = 32'h0;
    {bank3[1850], bank2[1850], bank1[1850], bank0[1850]} = 32'h0;
    {bank3[1851], bank2[1851], bank1[1851], bank0[1851]} = 32'h0;
    {bank3[1852], bank2[1852], bank1[1852], bank0[1852]} = 32'h0;
    {bank3[1853], bank2[1853], bank1[1853], bank0[1853]} = 32'h0;
    {bank3[1854], bank2[1854], bank1[1854], bank0[1854]} = 32'h0;
    {bank3[1855], bank2[1855], bank1[1855], bank0[1855]} = 32'h0;
    {bank3[1856], bank2[1856], bank1[1856], bank0[1856]} = 32'h0;
    {bank3[1857], bank2[1857], bank1[1857], bank0[1857]} = 32'h0;
    {bank3[1858], bank2[1858], bank1[1858], bank0[1858]} = 32'h0;
    {bank3[1859], bank2[1859], bank1[1859], bank0[1859]} = 32'h0;
    {bank3[1860], bank2[1860], bank1[1860], bank0[1860]} = 32'h0;
    {bank3[1861], bank2[1861], bank1[1861], bank0[1861]} = 32'h0;
    {bank3[1862], bank2[1862], bank1[1862], bank0[1862]} = 32'h0;
    {bank3[1863], bank2[1863], bank1[1863], bank0[1863]} = 32'h0;
    {bank3[1864], bank2[1864], bank1[1864], bank0[1864]} = 32'h0;
    {bank3[1865], bank2[1865], bank1[1865], bank0[1865]} = 32'h0;
    {bank3[1866], bank2[1866], bank1[1866], bank0[1866]} = 32'h0;
    {bank3[1867], bank2[1867], bank1[1867], bank0[1867]} = 32'h0;
    {bank3[1868], bank2[1868], bank1[1868], bank0[1868]} = 32'h0;
    {bank3[1869], bank2[1869], bank1[1869], bank0[1869]} = 32'h0;
    {bank3[1870], bank2[1870], bank1[1870], bank0[1870]} = 32'h0;
    {bank3[1871], bank2[1871], bank1[1871], bank0[1871]} = 32'h0;
    {bank3[1872], bank2[1872], bank1[1872], bank0[1872]} = 32'h0;
    {bank3[1873], bank2[1873], bank1[1873], bank0[1873]} = 32'h0;
    {bank3[1874], bank2[1874], bank1[1874], bank0[1874]} = 32'h0;
    {bank3[1875], bank2[1875], bank1[1875], bank0[1875]} = 32'h0;
    {bank3[1876], bank2[1876], bank1[1876], bank0[1876]} = 32'h0;
    {bank3[1877], bank2[1877], bank1[1877], bank0[1877]} = 32'h0;
    {bank3[1878], bank2[1878], bank1[1878], bank0[1878]} = 32'h0;
    {bank3[1879], bank2[1879], bank1[1879], bank0[1879]} = 32'h0;
    {bank3[1880], bank2[1880], bank1[1880], bank0[1880]} = 32'h0;
    {bank3[1881], bank2[1881], bank1[1881], bank0[1881]} = 32'h0;
    {bank3[1882], bank2[1882], bank1[1882], bank0[1882]} = 32'h0;
    {bank3[1883], bank2[1883], bank1[1883], bank0[1883]} = 32'h0;
    {bank3[1884], bank2[1884], bank1[1884], bank0[1884]} = 32'h0;
    {bank3[1885], bank2[1885], bank1[1885], bank0[1885]} = 32'h0;
    {bank3[1886], bank2[1886], bank1[1886], bank0[1886]} = 32'h0;
    {bank3[1887], bank2[1887], bank1[1887], bank0[1887]} = 32'h0;
    {bank3[1888], bank2[1888], bank1[1888], bank0[1888]} = 32'h0;
    {bank3[1889], bank2[1889], bank1[1889], bank0[1889]} = 32'h0;
    {bank3[1890], bank2[1890], bank1[1890], bank0[1890]} = 32'h0;
    {bank3[1891], bank2[1891], bank1[1891], bank0[1891]} = 32'h0;
    {bank3[1892], bank2[1892], bank1[1892], bank0[1892]} = 32'h0;
    {bank3[1893], bank2[1893], bank1[1893], bank0[1893]} = 32'h0;
    {bank3[1894], bank2[1894], bank1[1894], bank0[1894]} = 32'h0;
    {bank3[1895], bank2[1895], bank1[1895], bank0[1895]} = 32'h0;
    {bank3[1896], bank2[1896], bank1[1896], bank0[1896]} = 32'h0;
    {bank3[1897], bank2[1897], bank1[1897], bank0[1897]} = 32'h0;
    {bank3[1898], bank2[1898], bank1[1898], bank0[1898]} = 32'h0;
    {bank3[1899], bank2[1899], bank1[1899], bank0[1899]} = 32'h0;
    {bank3[1900], bank2[1900], bank1[1900], bank0[1900]} = 32'h0;
    {bank3[1901], bank2[1901], bank1[1901], bank0[1901]} = 32'h0;
    {bank3[1902], bank2[1902], bank1[1902], bank0[1902]} = 32'h0;
    {bank3[1903], bank2[1903], bank1[1903], bank0[1903]} = 32'h0;
    {bank3[1904], bank2[1904], bank1[1904], bank0[1904]} = 32'h0;
    {bank3[1905], bank2[1905], bank1[1905], bank0[1905]} = 32'h0;
    {bank3[1906], bank2[1906], bank1[1906], bank0[1906]} = 32'h0;
    {bank3[1907], bank2[1907], bank1[1907], bank0[1907]} = 32'h0;
    {bank3[1908], bank2[1908], bank1[1908], bank0[1908]} = 32'h0;
    {bank3[1909], bank2[1909], bank1[1909], bank0[1909]} = 32'h0;
    {bank3[1910], bank2[1910], bank1[1910], bank0[1910]} = 32'h0;
    {bank3[1911], bank2[1911], bank1[1911], bank0[1911]} = 32'h0;
    {bank3[1912], bank2[1912], bank1[1912], bank0[1912]} = 32'h0;
    {bank3[1913], bank2[1913], bank1[1913], bank0[1913]} = 32'h0;
    {bank3[1914], bank2[1914], bank1[1914], bank0[1914]} = 32'h0;
    {bank3[1915], bank2[1915], bank1[1915], bank0[1915]} = 32'h0;
    {bank3[1916], bank2[1916], bank1[1916], bank0[1916]} = 32'h0;
    {bank3[1917], bank2[1917], bank1[1917], bank0[1917]} = 32'h0;
    {bank3[1918], bank2[1918], bank1[1918], bank0[1918]} = 32'h0;
    {bank3[1919], bank2[1919], bank1[1919], bank0[1919]} = 32'h0;
    {bank3[1920], bank2[1920], bank1[1920], bank0[1920]} = 32'h0;
    {bank3[1921], bank2[1921], bank1[1921], bank0[1921]} = 32'h0;
    {bank3[1922], bank2[1922], bank1[1922], bank0[1922]} = 32'h0;
    {bank3[1923], bank2[1923], bank1[1923], bank0[1923]} = 32'h0;
    {bank3[1924], bank2[1924], bank1[1924], bank0[1924]} = 32'h0;
    {bank3[1925], bank2[1925], bank1[1925], bank0[1925]} = 32'h0;
    {bank3[1926], bank2[1926], bank1[1926], bank0[1926]} = 32'h0;
    {bank3[1927], bank2[1927], bank1[1927], bank0[1927]} = 32'h0;
    {bank3[1928], bank2[1928], bank1[1928], bank0[1928]} = 32'h0;
    {bank3[1929], bank2[1929], bank1[1929], bank0[1929]} = 32'h0;
    {bank3[1930], bank2[1930], bank1[1930], bank0[1930]} = 32'h0;
    {bank3[1931], bank2[1931], bank1[1931], bank0[1931]} = 32'h0;
    {bank3[1932], bank2[1932], bank1[1932], bank0[1932]} = 32'h0;
    {bank3[1933], bank2[1933], bank1[1933], bank0[1933]} = 32'h0;
    {bank3[1934], bank2[1934], bank1[1934], bank0[1934]} = 32'h0;
    {bank3[1935], bank2[1935], bank1[1935], bank0[1935]} = 32'h0;
    {bank3[1936], bank2[1936], bank1[1936], bank0[1936]} = 32'h0;
    {bank3[1937], bank2[1937], bank1[1937], bank0[1937]} = 32'h0;
    {bank3[1938], bank2[1938], bank1[1938], bank0[1938]} = 32'h0;
    {bank3[1939], bank2[1939], bank1[1939], bank0[1939]} = 32'h0;
    {bank3[1940], bank2[1940], bank1[1940], bank0[1940]} = 32'h0;
    {bank3[1941], bank2[1941], bank1[1941], bank0[1941]} = 32'h0;
    {bank3[1942], bank2[1942], bank1[1942], bank0[1942]} = 32'h0;
    {bank3[1943], bank2[1943], bank1[1943], bank0[1943]} = 32'h0;
    {bank3[1944], bank2[1944], bank1[1944], bank0[1944]} = 32'h0;
    {bank3[1945], bank2[1945], bank1[1945], bank0[1945]} = 32'h0;
    {bank3[1946], bank2[1946], bank1[1946], bank0[1946]} = 32'h0;
    {bank3[1947], bank2[1947], bank1[1947], bank0[1947]} = 32'h0;
    {bank3[1948], bank2[1948], bank1[1948], bank0[1948]} = 32'h0;
    {bank3[1949], bank2[1949], bank1[1949], bank0[1949]} = 32'h0;
    {bank3[1950], bank2[1950], bank1[1950], bank0[1950]} = 32'h0;
    {bank3[1951], bank2[1951], bank1[1951], bank0[1951]} = 32'h0;
    {bank3[1952], bank2[1952], bank1[1952], bank0[1952]} = 32'h0;
    {bank3[1953], bank2[1953], bank1[1953], bank0[1953]} = 32'h0;
    {bank3[1954], bank2[1954], bank1[1954], bank0[1954]} = 32'h0;
    {bank3[1955], bank2[1955], bank1[1955], bank0[1955]} = 32'h0;
    {bank3[1956], bank2[1956], bank1[1956], bank0[1956]} = 32'h0;
    {bank3[1957], bank2[1957], bank1[1957], bank0[1957]} = 32'h0;
    {bank3[1958], bank2[1958], bank1[1958], bank0[1958]} = 32'h0;
    {bank3[1959], bank2[1959], bank1[1959], bank0[1959]} = 32'h0;
    {bank3[1960], bank2[1960], bank1[1960], bank0[1960]} = 32'h0;
    {bank3[1961], bank2[1961], bank1[1961], bank0[1961]} = 32'h0;
    {bank3[1962], bank2[1962], bank1[1962], bank0[1962]} = 32'h0;
    {bank3[1963], bank2[1963], bank1[1963], bank0[1963]} = 32'h0;
    {bank3[1964], bank2[1964], bank1[1964], bank0[1964]} = 32'h0;
    {bank3[1965], bank2[1965], bank1[1965], bank0[1965]} = 32'h0;
    {bank3[1966], bank2[1966], bank1[1966], bank0[1966]} = 32'h0;
    {bank3[1967], bank2[1967], bank1[1967], bank0[1967]} = 32'h0;
    {bank3[1968], bank2[1968], bank1[1968], bank0[1968]} = 32'h0;
    {bank3[1969], bank2[1969], bank1[1969], bank0[1969]} = 32'h0;
    {bank3[1970], bank2[1970], bank1[1970], bank0[1970]} = 32'h0;
    {bank3[1971], bank2[1971], bank1[1971], bank0[1971]} = 32'h0;
    {bank3[1972], bank2[1972], bank1[1972], bank0[1972]} = 32'h0;
    {bank3[1973], bank2[1973], bank1[1973], bank0[1973]} = 32'h0;
    {bank3[1974], bank2[1974], bank1[1974], bank0[1974]} = 32'h0;
    {bank3[1975], bank2[1975], bank1[1975], bank0[1975]} = 32'h0;
    {bank3[1976], bank2[1976], bank1[1976], bank0[1976]} = 32'h0;
    {bank3[1977], bank2[1977], bank1[1977], bank0[1977]} = 32'h0;
    {bank3[1978], bank2[1978], bank1[1978], bank0[1978]} = 32'h0;
    {bank3[1979], bank2[1979], bank1[1979], bank0[1979]} = 32'h0;
    {bank3[1980], bank2[1980], bank1[1980], bank0[1980]} = 32'h0;
    {bank3[1981], bank2[1981], bank1[1981], bank0[1981]} = 32'h0;
    {bank3[1982], bank2[1982], bank1[1982], bank0[1982]} = 32'h0;
    {bank3[1983], bank2[1983], bank1[1983], bank0[1983]} = 32'h0;
    {bank3[1984], bank2[1984], bank1[1984], bank0[1984]} = 32'h0;
    {bank3[1985], bank2[1985], bank1[1985], bank0[1985]} = 32'h0;
    {bank3[1986], bank2[1986], bank1[1986], bank0[1986]} = 32'h0;
    {bank3[1987], bank2[1987], bank1[1987], bank0[1987]} = 32'h0;
    {bank3[1988], bank2[1988], bank1[1988], bank0[1988]} = 32'h0;
    {bank3[1989], bank2[1989], bank1[1989], bank0[1989]} = 32'h0;
    {bank3[1990], bank2[1990], bank1[1990], bank0[1990]} = 32'h0;
    {bank3[1991], bank2[1991], bank1[1991], bank0[1991]} = 32'h0;
    {bank3[1992], bank2[1992], bank1[1992], bank0[1992]} = 32'h0;
    {bank3[1993], bank2[1993], bank1[1993], bank0[1993]} = 32'h0;
    {bank3[1994], bank2[1994], bank1[1994], bank0[1994]} = 32'h0;
    {bank3[1995], bank2[1995], bank1[1995], bank0[1995]} = 32'h0;
    {bank3[1996], bank2[1996], bank1[1996], bank0[1996]} = 32'h0;
    {bank3[1997], bank2[1997], bank1[1997], bank0[1997]} = 32'h0;
    {bank3[1998], bank2[1998], bank1[1998], bank0[1998]} = 32'h0;
    {bank3[1999], bank2[1999], bank1[1999], bank0[1999]} = 32'h0;
    {bank3[2000], bank2[2000], bank1[2000], bank0[2000]} = 32'h0;
    {bank3[2001], bank2[2001], bank1[2001], bank0[2001]} = 32'h0;
    {bank3[2002], bank2[2002], bank1[2002], bank0[2002]} = 32'h0;
    {bank3[2003], bank2[2003], bank1[2003], bank0[2003]} = 32'h0;
    {bank3[2004], bank2[2004], bank1[2004], bank0[2004]} = 32'h0;
    {bank3[2005], bank2[2005], bank1[2005], bank0[2005]} = 32'h0;
    {bank3[2006], bank2[2006], bank1[2006], bank0[2006]} = 32'h0;
    {bank3[2007], bank2[2007], bank1[2007], bank0[2007]} = 32'h0;
    {bank3[2008], bank2[2008], bank1[2008], bank0[2008]} = 32'h0;
    {bank3[2009], bank2[2009], bank1[2009], bank0[2009]} = 32'h0;
    {bank3[2010], bank2[2010], bank1[2010], bank0[2010]} = 32'h0;
    {bank3[2011], bank2[2011], bank1[2011], bank0[2011]} = 32'h0;
    {bank3[2012], bank2[2012], bank1[2012], bank0[2012]} = 32'h0;
    {bank3[2013], bank2[2013], bank1[2013], bank0[2013]} = 32'h0;
    {bank3[2014], bank2[2014], bank1[2014], bank0[2014]} = 32'h0;
    {bank3[2015], bank2[2015], bank1[2015], bank0[2015]} = 32'h0;
    {bank3[2016], bank2[2016], bank1[2016], bank0[2016]} = 32'h0;
    {bank3[2017], bank2[2017], bank1[2017], bank0[2017]} = 32'h0;
    {bank3[2018], bank2[2018], bank1[2018], bank0[2018]} = 32'h0;
    {bank3[2019], bank2[2019], bank1[2019], bank0[2019]} = 32'h0;
    {bank3[2020], bank2[2020], bank1[2020], bank0[2020]} = 32'h0;
    {bank3[2021], bank2[2021], bank1[2021], bank0[2021]} = 32'h0;
    {bank3[2022], bank2[2022], bank1[2022], bank0[2022]} = 32'h0;
    {bank3[2023], bank2[2023], bank1[2023], bank0[2023]} = 32'h0;
    {bank3[2024], bank2[2024], bank1[2024], bank0[2024]} = 32'h0;
    {bank3[2025], bank2[2025], bank1[2025], bank0[2025]} = 32'h0;
    {bank3[2026], bank2[2026], bank1[2026], bank0[2026]} = 32'h0;
    {bank3[2027], bank2[2027], bank1[2027], bank0[2027]} = 32'h0;
    {bank3[2028], bank2[2028], bank1[2028], bank0[2028]} = 32'h0;
    {bank3[2029], bank2[2029], bank1[2029], bank0[2029]} = 32'h0;
    {bank3[2030], bank2[2030], bank1[2030], bank0[2030]} = 32'h0;
    {bank3[2031], bank2[2031], bank1[2031], bank0[2031]} = 32'h0;
    {bank3[2032], bank2[2032], bank1[2032], bank0[2032]} = 32'h0;
    {bank3[2033], bank2[2033], bank1[2033], bank0[2033]} = 32'h0;
    {bank3[2034], bank2[2034], bank1[2034], bank0[2034]} = 32'h0;
    {bank3[2035], bank2[2035], bank1[2035], bank0[2035]} = 32'h0;
    {bank3[2036], bank2[2036], bank1[2036], bank0[2036]} = 32'h0;
    {bank3[2037], bank2[2037], bank1[2037], bank0[2037]} = 32'h0;
    {bank3[2038], bank2[2038], bank1[2038], bank0[2038]} = 32'h0;
    {bank3[2039], bank2[2039], bank1[2039], bank0[2039]} = 32'h0;
    {bank3[2040], bank2[2040], bank1[2040], bank0[2040]} = 32'h0;
    {bank3[2041], bank2[2041], bank1[2041], bank0[2041]} = 32'h0;
    {bank3[2042], bank2[2042], bank1[2042], bank0[2042]} = 32'h0;
    {bank3[2043], bank2[2043], bank1[2043], bank0[2043]} = 32'h0;
    {bank3[2044], bank2[2044], bank1[2044], bank0[2044]} = 32'h0;
    {bank3[2045], bank2[2045], bank1[2045], bank0[2045]} = 32'h0;
    {bank3[2046], bank2[2046], bank1[2046], bank0[2046]} = 32'h0;
    {bank3[2047], bank2[2047], bank1[2047], bank0[2047]} = 32'h0;
    {bank3[2048], bank2[2048], bank1[2048], bank0[2048]} = 32'h0;
    {bank3[2049], bank2[2049], bank1[2049], bank0[2049]} = 32'h0;
    {bank3[2050], bank2[2050], bank1[2050], bank0[2050]} = 32'h0;
    {bank3[2051], bank2[2051], bank1[2051], bank0[2051]} = 32'h0;
    {bank3[2052], bank2[2052], bank1[2052], bank0[2052]} = 32'h0;
    {bank3[2053], bank2[2053], bank1[2053], bank0[2053]} = 32'h0;
    {bank3[2054], bank2[2054], bank1[2054], bank0[2054]} = 32'h0;
    {bank3[2055], bank2[2055], bank1[2055], bank0[2055]} = 32'h0;
    {bank3[2056], bank2[2056], bank1[2056], bank0[2056]} = 32'h0;
    {bank3[2057], bank2[2057], bank1[2057], bank0[2057]} = 32'h0;
    {bank3[2058], bank2[2058], bank1[2058], bank0[2058]} = 32'h0;
    {bank3[2059], bank2[2059], bank1[2059], bank0[2059]} = 32'h0;
    {bank3[2060], bank2[2060], bank1[2060], bank0[2060]} = 32'h0;
    {bank3[2061], bank2[2061], bank1[2061], bank0[2061]} = 32'h0;
    {bank3[2062], bank2[2062], bank1[2062], bank0[2062]} = 32'h0;
    {bank3[2063], bank2[2063], bank1[2063], bank0[2063]} = 32'h0;
    {bank3[2064], bank2[2064], bank1[2064], bank0[2064]} = 32'h0;
    {bank3[2065], bank2[2065], bank1[2065], bank0[2065]} = 32'h0;
    {bank3[2066], bank2[2066], bank1[2066], bank0[2066]} = 32'h0;
    {bank3[2067], bank2[2067], bank1[2067], bank0[2067]} = 32'h0;
    {bank3[2068], bank2[2068], bank1[2068], bank0[2068]} = 32'h0;
    {bank3[2069], bank2[2069], bank1[2069], bank0[2069]} = 32'h0;
    {bank3[2070], bank2[2070], bank1[2070], bank0[2070]} = 32'h0;
    {bank3[2071], bank2[2071], bank1[2071], bank0[2071]} = 32'h0;
    {bank3[2072], bank2[2072], bank1[2072], bank0[2072]} = 32'h0;
    {bank3[2073], bank2[2073], bank1[2073], bank0[2073]} = 32'h0;
    {bank3[2074], bank2[2074], bank1[2074], bank0[2074]} = 32'h0;
    {bank3[2075], bank2[2075], bank1[2075], bank0[2075]} = 32'h0;
    {bank3[2076], bank2[2076], bank1[2076], bank0[2076]} = 32'h0;
    {bank3[2077], bank2[2077], bank1[2077], bank0[2077]} = 32'h0;
    {bank3[2078], bank2[2078], bank1[2078], bank0[2078]} = 32'h0;
    {bank3[2079], bank2[2079], bank1[2079], bank0[2079]} = 32'h0;
    {bank3[2080], bank2[2080], bank1[2080], bank0[2080]} = 32'h0;
    {bank3[2081], bank2[2081], bank1[2081], bank0[2081]} = 32'h0;
    {bank3[2082], bank2[2082], bank1[2082], bank0[2082]} = 32'h0;
    {bank3[2083], bank2[2083], bank1[2083], bank0[2083]} = 32'h0;
    {bank3[2084], bank2[2084], bank1[2084], bank0[2084]} = 32'h0;
    {bank3[2085], bank2[2085], bank1[2085], bank0[2085]} = 32'h0;
    {bank3[2086], bank2[2086], bank1[2086], bank0[2086]} = 32'h0;
    {bank3[2087], bank2[2087], bank1[2087], bank0[2087]} = 32'h0;
    {bank3[2088], bank2[2088], bank1[2088], bank0[2088]} = 32'h0;
    {bank3[2089], bank2[2089], bank1[2089], bank0[2089]} = 32'h0;
    {bank3[2090], bank2[2090], bank1[2090], bank0[2090]} = 32'h0;
    {bank3[2091], bank2[2091], bank1[2091], bank0[2091]} = 32'h0;
    {bank3[2092], bank2[2092], bank1[2092], bank0[2092]} = 32'h0;
    {bank3[2093], bank2[2093], bank1[2093], bank0[2093]} = 32'h0;
    {bank3[2094], bank2[2094], bank1[2094], bank0[2094]} = 32'h0;
    {bank3[2095], bank2[2095], bank1[2095], bank0[2095]} = 32'h0;
    {bank3[2096], bank2[2096], bank1[2096], bank0[2096]} = 32'h0;
    {bank3[2097], bank2[2097], bank1[2097], bank0[2097]} = 32'h0;
    {bank3[2098], bank2[2098], bank1[2098], bank0[2098]} = 32'h0;
    {bank3[2099], bank2[2099], bank1[2099], bank0[2099]} = 32'h0;
    {bank3[2100], bank2[2100], bank1[2100], bank0[2100]} = 32'h0;
    {bank3[2101], bank2[2101], bank1[2101], bank0[2101]} = 32'h0;
    {bank3[2102], bank2[2102], bank1[2102], bank0[2102]} = 32'h0;
    {bank3[2103], bank2[2103], bank1[2103], bank0[2103]} = 32'h0;
    {bank3[2104], bank2[2104], bank1[2104], bank0[2104]} = 32'h0;
    {bank3[2105], bank2[2105], bank1[2105], bank0[2105]} = 32'h0;
    {bank3[2106], bank2[2106], bank1[2106], bank0[2106]} = 32'h0;
    {bank3[2107], bank2[2107], bank1[2107], bank0[2107]} = 32'h0;
    {bank3[2108], bank2[2108], bank1[2108], bank0[2108]} = 32'h0;
    {bank3[2109], bank2[2109], bank1[2109], bank0[2109]} = 32'h0;
    {bank3[2110], bank2[2110], bank1[2110], bank0[2110]} = 32'h0;
    {bank3[2111], bank2[2111], bank1[2111], bank0[2111]} = 32'h0;
    {bank3[2112], bank2[2112], bank1[2112], bank0[2112]} = 32'h0;
    {bank3[2113], bank2[2113], bank1[2113], bank0[2113]} = 32'h0;
    {bank3[2114], bank2[2114], bank1[2114], bank0[2114]} = 32'h0;
    {bank3[2115], bank2[2115], bank1[2115], bank0[2115]} = 32'h0;
    {bank3[2116], bank2[2116], bank1[2116], bank0[2116]} = 32'h0;
    {bank3[2117], bank2[2117], bank1[2117], bank0[2117]} = 32'h0;
    {bank3[2118], bank2[2118], bank1[2118], bank0[2118]} = 32'h0;
    {bank3[2119], bank2[2119], bank1[2119], bank0[2119]} = 32'h0;
    {bank3[2120], bank2[2120], bank1[2120], bank0[2120]} = 32'h0;
    {bank3[2121], bank2[2121], bank1[2121], bank0[2121]} = 32'h0;
    {bank3[2122], bank2[2122], bank1[2122], bank0[2122]} = 32'h0;
    {bank3[2123], bank2[2123], bank1[2123], bank0[2123]} = 32'h0;
    {bank3[2124], bank2[2124], bank1[2124], bank0[2124]} = 32'h0;
    {bank3[2125], bank2[2125], bank1[2125], bank0[2125]} = 32'h0;
    {bank3[2126], bank2[2126], bank1[2126], bank0[2126]} = 32'h0;
    {bank3[2127], bank2[2127], bank1[2127], bank0[2127]} = 32'h0;
    {bank3[2128], bank2[2128], bank1[2128], bank0[2128]} = 32'h0;
    {bank3[2129], bank2[2129], bank1[2129], bank0[2129]} = 32'h0;
    {bank3[2130], bank2[2130], bank1[2130], bank0[2130]} = 32'h0;
    {bank3[2131], bank2[2131], bank1[2131], bank0[2131]} = 32'h0;
    {bank3[2132], bank2[2132], bank1[2132], bank0[2132]} = 32'h0;
    {bank3[2133], bank2[2133], bank1[2133], bank0[2133]} = 32'h0;
    {bank3[2134], bank2[2134], bank1[2134], bank0[2134]} = 32'h0;
    {bank3[2135], bank2[2135], bank1[2135], bank0[2135]} = 32'h0;
    {bank3[2136], bank2[2136], bank1[2136], bank0[2136]} = 32'h0;
    {bank3[2137], bank2[2137], bank1[2137], bank0[2137]} = 32'h0;
    {bank3[2138], bank2[2138], bank1[2138], bank0[2138]} = 32'h0;
    {bank3[2139], bank2[2139], bank1[2139], bank0[2139]} = 32'h0;
    {bank3[2140], bank2[2140], bank1[2140], bank0[2140]} = 32'h0;
    {bank3[2141], bank2[2141], bank1[2141], bank0[2141]} = 32'h0;
    {bank3[2142], bank2[2142], bank1[2142], bank0[2142]} = 32'h0;
    {bank3[2143], bank2[2143], bank1[2143], bank0[2143]} = 32'h0;
    {bank3[2144], bank2[2144], bank1[2144], bank0[2144]} = 32'h0;
    {bank3[2145], bank2[2145], bank1[2145], bank0[2145]} = 32'h0;
    {bank3[2146], bank2[2146], bank1[2146], bank0[2146]} = 32'h0;
    {bank3[2147], bank2[2147], bank1[2147], bank0[2147]} = 32'h0;
    {bank3[2148], bank2[2148], bank1[2148], bank0[2148]} = 32'h0;
    {bank3[2149], bank2[2149], bank1[2149], bank0[2149]} = 32'h0;
    {bank3[2150], bank2[2150], bank1[2150], bank0[2150]} = 32'h0;
    {bank3[2151], bank2[2151], bank1[2151], bank0[2151]} = 32'h0;
    {bank3[2152], bank2[2152], bank1[2152], bank0[2152]} = 32'h0;
    {bank3[2153], bank2[2153], bank1[2153], bank0[2153]} = 32'h0;
    {bank3[2154], bank2[2154], bank1[2154], bank0[2154]} = 32'h0;
    {bank3[2155], bank2[2155], bank1[2155], bank0[2155]} = 32'h0;
    {bank3[2156], bank2[2156], bank1[2156], bank0[2156]} = 32'h0;
    {bank3[2157], bank2[2157], bank1[2157], bank0[2157]} = 32'h0;
    {bank3[2158], bank2[2158], bank1[2158], bank0[2158]} = 32'h0;
    {bank3[2159], bank2[2159], bank1[2159], bank0[2159]} = 32'h0;
    {bank3[2160], bank2[2160], bank1[2160], bank0[2160]} = 32'h0;
    {bank3[2161], bank2[2161], bank1[2161], bank0[2161]} = 32'h0;
    {bank3[2162], bank2[2162], bank1[2162], bank0[2162]} = 32'h0;
    {bank3[2163], bank2[2163], bank1[2163], bank0[2163]} = 32'h0;
    {bank3[2164], bank2[2164], bank1[2164], bank0[2164]} = 32'h0;
    {bank3[2165], bank2[2165], bank1[2165], bank0[2165]} = 32'h0;
    {bank3[2166], bank2[2166], bank1[2166], bank0[2166]} = 32'h0;
    {bank3[2167], bank2[2167], bank1[2167], bank0[2167]} = 32'h0;
    {bank3[2168], bank2[2168], bank1[2168], bank0[2168]} = 32'h0;
    {bank3[2169], bank2[2169], bank1[2169], bank0[2169]} = 32'h0;
    {bank3[2170], bank2[2170], bank1[2170], bank0[2170]} = 32'h0;
    {bank3[2171], bank2[2171], bank1[2171], bank0[2171]} = 32'h0;
    {bank3[2172], bank2[2172], bank1[2172], bank0[2172]} = 32'h0;
    {bank3[2173], bank2[2173], bank1[2173], bank0[2173]} = 32'h0;
    {bank3[2174], bank2[2174], bank1[2174], bank0[2174]} = 32'h0;
    {bank3[2175], bank2[2175], bank1[2175], bank0[2175]} = 32'h0;
    {bank3[2176], bank2[2176], bank1[2176], bank0[2176]} = 32'h0;
    {bank3[2177], bank2[2177], bank1[2177], bank0[2177]} = 32'h0;
    {bank3[2178], bank2[2178], bank1[2178], bank0[2178]} = 32'h0;
    {bank3[2179], bank2[2179], bank1[2179], bank0[2179]} = 32'h0;
    {bank3[2180], bank2[2180], bank1[2180], bank0[2180]} = 32'h0;
    {bank3[2181], bank2[2181], bank1[2181], bank0[2181]} = 32'h0;
    {bank3[2182], bank2[2182], bank1[2182], bank0[2182]} = 32'h0;
    {bank3[2183], bank2[2183], bank1[2183], bank0[2183]} = 32'h0;
    {bank3[2184], bank2[2184], bank1[2184], bank0[2184]} = 32'h0;
    {bank3[2185], bank2[2185], bank1[2185], bank0[2185]} = 32'h0;
    {bank3[2186], bank2[2186], bank1[2186], bank0[2186]} = 32'h0;
    {bank3[2187], bank2[2187], bank1[2187], bank0[2187]} = 32'h0;
    {bank3[2188], bank2[2188], bank1[2188], bank0[2188]} = 32'h0;
    {bank3[2189], bank2[2189], bank1[2189], bank0[2189]} = 32'h0;
    {bank3[2190], bank2[2190], bank1[2190], bank0[2190]} = 32'h0;
    {bank3[2191], bank2[2191], bank1[2191], bank0[2191]} = 32'h0;
    {bank3[2192], bank2[2192], bank1[2192], bank0[2192]} = 32'h0;
    {bank3[2193], bank2[2193], bank1[2193], bank0[2193]} = 32'h0;
    {bank3[2194], bank2[2194], bank1[2194], bank0[2194]} = 32'h0;
    {bank3[2195], bank2[2195], bank1[2195], bank0[2195]} = 32'h0;
    {bank3[2196], bank2[2196], bank1[2196], bank0[2196]} = 32'h0;
    {bank3[2197], bank2[2197], bank1[2197], bank0[2197]} = 32'h0;
    {bank3[2198], bank2[2198], bank1[2198], bank0[2198]} = 32'h0;
    {bank3[2199], bank2[2199], bank1[2199], bank0[2199]} = 32'h0;
    {bank3[2200], bank2[2200], bank1[2200], bank0[2200]} = 32'h0;
    {bank3[2201], bank2[2201], bank1[2201], bank0[2201]} = 32'h0;
    {bank3[2202], bank2[2202], bank1[2202], bank0[2202]} = 32'h0;
    {bank3[2203], bank2[2203], bank1[2203], bank0[2203]} = 32'h0;
    {bank3[2204], bank2[2204], bank1[2204], bank0[2204]} = 32'h0;
    {bank3[2205], bank2[2205], bank1[2205], bank0[2205]} = 32'h0;
    {bank3[2206], bank2[2206], bank1[2206], bank0[2206]} = 32'h0;
    {bank3[2207], bank2[2207], bank1[2207], bank0[2207]} = 32'h0;
    {bank3[2208], bank2[2208], bank1[2208], bank0[2208]} = 32'h0;
    {bank3[2209], bank2[2209], bank1[2209], bank0[2209]} = 32'h0;
    {bank3[2210], bank2[2210], bank1[2210], bank0[2210]} = 32'h0;
    {bank3[2211], bank2[2211], bank1[2211], bank0[2211]} = 32'h0;
    {bank3[2212], bank2[2212], bank1[2212], bank0[2212]} = 32'h0;
    {bank3[2213], bank2[2213], bank1[2213], bank0[2213]} = 32'h0;
    {bank3[2214], bank2[2214], bank1[2214], bank0[2214]} = 32'h0;
    {bank3[2215], bank2[2215], bank1[2215], bank0[2215]} = 32'h0;
    {bank3[2216], bank2[2216], bank1[2216], bank0[2216]} = 32'h0;
    {bank3[2217], bank2[2217], bank1[2217], bank0[2217]} = 32'h0;
    {bank3[2218], bank2[2218], bank1[2218], bank0[2218]} = 32'h0;
    {bank3[2219], bank2[2219], bank1[2219], bank0[2219]} = 32'h0;
    {bank3[2220], bank2[2220], bank1[2220], bank0[2220]} = 32'h0;
    {bank3[2221], bank2[2221], bank1[2221], bank0[2221]} = 32'h0;
    {bank3[2222], bank2[2222], bank1[2222], bank0[2222]} = 32'h0;
    {bank3[2223], bank2[2223], bank1[2223], bank0[2223]} = 32'h0;
    {bank3[2224], bank2[2224], bank1[2224], bank0[2224]} = 32'h0;
    {bank3[2225], bank2[2225], bank1[2225], bank0[2225]} = 32'h0;
    {bank3[2226], bank2[2226], bank1[2226], bank0[2226]} = 32'h0;
    {bank3[2227], bank2[2227], bank1[2227], bank0[2227]} = 32'h0;
    {bank3[2228], bank2[2228], bank1[2228], bank0[2228]} = 32'h0;
    {bank3[2229], bank2[2229], bank1[2229], bank0[2229]} = 32'h0;
    {bank3[2230], bank2[2230], bank1[2230], bank0[2230]} = 32'h0;
    {bank3[2231], bank2[2231], bank1[2231], bank0[2231]} = 32'h0;
    {bank3[2232], bank2[2232], bank1[2232], bank0[2232]} = 32'h0;
    {bank3[2233], bank2[2233], bank1[2233], bank0[2233]} = 32'h0;
    {bank3[2234], bank2[2234], bank1[2234], bank0[2234]} = 32'h0;
    {bank3[2235], bank2[2235], bank1[2235], bank0[2235]} = 32'h0;
    {bank3[2236], bank2[2236], bank1[2236], bank0[2236]} = 32'h0;
    {bank3[2237], bank2[2237], bank1[2237], bank0[2237]} = 32'h0;
    {bank3[2238], bank2[2238], bank1[2238], bank0[2238]} = 32'h0;
    {bank3[2239], bank2[2239], bank1[2239], bank0[2239]} = 32'h0;
    {bank3[2240], bank2[2240], bank1[2240], bank0[2240]} = 32'h0;
    {bank3[2241], bank2[2241], bank1[2241], bank0[2241]} = 32'h0;
    {bank3[2242], bank2[2242], bank1[2242], bank0[2242]} = 32'h0;
    {bank3[2243], bank2[2243], bank1[2243], bank0[2243]} = 32'h0;
    {bank3[2244], bank2[2244], bank1[2244], bank0[2244]} = 32'h0;
    {bank3[2245], bank2[2245], bank1[2245], bank0[2245]} = 32'h0;
    {bank3[2246], bank2[2246], bank1[2246], bank0[2246]} = 32'h0;
    {bank3[2247], bank2[2247], bank1[2247], bank0[2247]} = 32'h0;
    {bank3[2248], bank2[2248], bank1[2248], bank0[2248]} = 32'h0;
    {bank3[2249], bank2[2249], bank1[2249], bank0[2249]} = 32'h0;
    {bank3[2250], bank2[2250], bank1[2250], bank0[2250]} = 32'h0;
    {bank3[2251], bank2[2251], bank1[2251], bank0[2251]} = 32'h0;
    {bank3[2252], bank2[2252], bank1[2252], bank0[2252]} = 32'h0;
    {bank3[2253], bank2[2253], bank1[2253], bank0[2253]} = 32'h0;
    {bank3[2254], bank2[2254], bank1[2254], bank0[2254]} = 32'h0;
    {bank3[2255], bank2[2255], bank1[2255], bank0[2255]} = 32'h0;
    {bank3[2256], bank2[2256], bank1[2256], bank0[2256]} = 32'h0;
    {bank3[2257], bank2[2257], bank1[2257], bank0[2257]} = 32'h0;
    {bank3[2258], bank2[2258], bank1[2258], bank0[2258]} = 32'h0;
    {bank3[2259], bank2[2259], bank1[2259], bank0[2259]} = 32'h0;
    {bank3[2260], bank2[2260], bank1[2260], bank0[2260]} = 32'h0;
    {bank3[2261], bank2[2261], bank1[2261], bank0[2261]} = 32'h0;
    {bank3[2262], bank2[2262], bank1[2262], bank0[2262]} = 32'h0;
    {bank3[2263], bank2[2263], bank1[2263], bank0[2263]} = 32'h0;
    {bank3[2264], bank2[2264], bank1[2264], bank0[2264]} = 32'h0;
    {bank3[2265], bank2[2265], bank1[2265], bank0[2265]} = 32'h0;
    {bank3[2266], bank2[2266], bank1[2266], bank0[2266]} = 32'h0;
    {bank3[2267], bank2[2267], bank1[2267], bank0[2267]} = 32'h0;
    {bank3[2268], bank2[2268], bank1[2268], bank0[2268]} = 32'h0;
    {bank3[2269], bank2[2269], bank1[2269], bank0[2269]} = 32'h0;
    {bank3[2270], bank2[2270], bank1[2270], bank0[2270]} = 32'h0;
    {bank3[2271], bank2[2271], bank1[2271], bank0[2271]} = 32'h0;
    {bank3[2272], bank2[2272], bank1[2272], bank0[2272]} = 32'h0;
    {bank3[2273], bank2[2273], bank1[2273], bank0[2273]} = 32'h0;
    {bank3[2274], bank2[2274], bank1[2274], bank0[2274]} = 32'h0;
    {bank3[2275], bank2[2275], bank1[2275], bank0[2275]} = 32'h0;
    {bank3[2276], bank2[2276], bank1[2276], bank0[2276]} = 32'h0;
    {bank3[2277], bank2[2277], bank1[2277], bank0[2277]} = 32'h0;
    {bank3[2278], bank2[2278], bank1[2278], bank0[2278]} = 32'h0;
    {bank3[2279], bank2[2279], bank1[2279], bank0[2279]} = 32'h0;
    {bank3[2280], bank2[2280], bank1[2280], bank0[2280]} = 32'h0;
    {bank3[2281], bank2[2281], bank1[2281], bank0[2281]} = 32'h0;
    {bank3[2282], bank2[2282], bank1[2282], bank0[2282]} = 32'h0;
    {bank3[2283], bank2[2283], bank1[2283], bank0[2283]} = 32'h0;
    {bank3[2284], bank2[2284], bank1[2284], bank0[2284]} = 32'h0;
    {bank3[2285], bank2[2285], bank1[2285], bank0[2285]} = 32'h0;
    {bank3[2286], bank2[2286], bank1[2286], bank0[2286]} = 32'h0;
    {bank3[2287], bank2[2287], bank1[2287], bank0[2287]} = 32'h0;
    {bank3[2288], bank2[2288], bank1[2288], bank0[2288]} = 32'h0;
    {bank3[2289], bank2[2289], bank1[2289], bank0[2289]} = 32'h0;
    {bank3[2290], bank2[2290], bank1[2290], bank0[2290]} = 32'h0;
    {bank3[2291], bank2[2291], bank1[2291], bank0[2291]} = 32'h0;
    {bank3[2292], bank2[2292], bank1[2292], bank0[2292]} = 32'h0;
    {bank3[2293], bank2[2293], bank1[2293], bank0[2293]} = 32'h0;
    {bank3[2294], bank2[2294], bank1[2294], bank0[2294]} = 32'h0;
    {bank3[2295], bank2[2295], bank1[2295], bank0[2295]} = 32'h0;
    {bank3[2296], bank2[2296], bank1[2296], bank0[2296]} = 32'h0;
    {bank3[2297], bank2[2297], bank1[2297], bank0[2297]} = 32'h0;
    {bank3[2298], bank2[2298], bank1[2298], bank0[2298]} = 32'h0;
    {bank3[2299], bank2[2299], bank1[2299], bank0[2299]} = 32'h0;
    {bank3[2300], bank2[2300], bank1[2300], bank0[2300]} = 32'h0;
    {bank3[2301], bank2[2301], bank1[2301], bank0[2301]} = 32'h0;
    {bank3[2302], bank2[2302], bank1[2302], bank0[2302]} = 32'h0;
    {bank3[2303], bank2[2303], bank1[2303], bank0[2303]} = 32'h0;
    {bank3[2304], bank2[2304], bank1[2304], bank0[2304]} = 32'h0;
    {bank3[2305], bank2[2305], bank1[2305], bank0[2305]} = 32'h0;
    {bank3[2306], bank2[2306], bank1[2306], bank0[2306]} = 32'h0;
    {bank3[2307], bank2[2307], bank1[2307], bank0[2307]} = 32'h0;
    {bank3[2308], bank2[2308], bank1[2308], bank0[2308]} = 32'h0;
    {bank3[2309], bank2[2309], bank1[2309], bank0[2309]} = 32'h0;
    {bank3[2310], bank2[2310], bank1[2310], bank0[2310]} = 32'h0;
    {bank3[2311], bank2[2311], bank1[2311], bank0[2311]} = 32'h0;
    {bank3[2312], bank2[2312], bank1[2312], bank0[2312]} = 32'h0;
    {bank3[2313], bank2[2313], bank1[2313], bank0[2313]} = 32'h0;
    {bank3[2314], bank2[2314], bank1[2314], bank0[2314]} = 32'h0;
    {bank3[2315], bank2[2315], bank1[2315], bank0[2315]} = 32'h0;
    {bank3[2316], bank2[2316], bank1[2316], bank0[2316]} = 32'h0;
    {bank3[2317], bank2[2317], bank1[2317], bank0[2317]} = 32'h0;
    {bank3[2318], bank2[2318], bank1[2318], bank0[2318]} = 32'h0;
    {bank3[2319], bank2[2319], bank1[2319], bank0[2319]} = 32'h0;
    {bank3[2320], bank2[2320], bank1[2320], bank0[2320]} = 32'h0;
    {bank3[2321], bank2[2321], bank1[2321], bank0[2321]} = 32'h0;
    {bank3[2322], bank2[2322], bank1[2322], bank0[2322]} = 32'h0;
    {bank3[2323], bank2[2323], bank1[2323], bank0[2323]} = 32'h0;
    {bank3[2324], bank2[2324], bank1[2324], bank0[2324]} = 32'h0;
    {bank3[2325], bank2[2325], bank1[2325], bank0[2325]} = 32'h0;
    {bank3[2326], bank2[2326], bank1[2326], bank0[2326]} = 32'h0;
    {bank3[2327], bank2[2327], bank1[2327], bank0[2327]} = 32'h0;
    {bank3[2328], bank2[2328], bank1[2328], bank0[2328]} = 32'h0;
    {bank3[2329], bank2[2329], bank1[2329], bank0[2329]} = 32'h0;
    {bank3[2330], bank2[2330], bank1[2330], bank0[2330]} = 32'h0;
    {bank3[2331], bank2[2331], bank1[2331], bank0[2331]} = 32'h0;
    {bank3[2332], bank2[2332], bank1[2332], bank0[2332]} = 32'h0;
    {bank3[2333], bank2[2333], bank1[2333], bank0[2333]} = 32'h0;
    {bank3[2334], bank2[2334], bank1[2334], bank0[2334]} = 32'h0;
    {bank3[2335], bank2[2335], bank1[2335], bank0[2335]} = 32'h0;
    {bank3[2336], bank2[2336], bank1[2336], bank0[2336]} = 32'h0;
    {bank3[2337], bank2[2337], bank1[2337], bank0[2337]} = 32'h0;
    {bank3[2338], bank2[2338], bank1[2338], bank0[2338]} = 32'h0;
    {bank3[2339], bank2[2339], bank1[2339], bank0[2339]} = 32'h0;
    {bank3[2340], bank2[2340], bank1[2340], bank0[2340]} = 32'h0;
    {bank3[2341], bank2[2341], bank1[2341], bank0[2341]} = 32'h0;
    {bank3[2342], bank2[2342], bank1[2342], bank0[2342]} = 32'h0;
    {bank3[2343], bank2[2343], bank1[2343], bank0[2343]} = 32'h0;
    {bank3[2344], bank2[2344], bank1[2344], bank0[2344]} = 32'h0;
    {bank3[2345], bank2[2345], bank1[2345], bank0[2345]} = 32'h0;
    {bank3[2346], bank2[2346], bank1[2346], bank0[2346]} = 32'h0;
    {bank3[2347], bank2[2347], bank1[2347], bank0[2347]} = 32'h0;
    {bank3[2348], bank2[2348], bank1[2348], bank0[2348]} = 32'h0;
    {bank3[2349], bank2[2349], bank1[2349], bank0[2349]} = 32'h0;
    {bank3[2350], bank2[2350], bank1[2350], bank0[2350]} = 32'h0;
    {bank3[2351], bank2[2351], bank1[2351], bank0[2351]} = 32'h0;
    {bank3[2352], bank2[2352], bank1[2352], bank0[2352]} = 32'h0;
    {bank3[2353], bank2[2353], bank1[2353], bank0[2353]} = 32'h0;
    {bank3[2354], bank2[2354], bank1[2354], bank0[2354]} = 32'h0;
    {bank3[2355], bank2[2355], bank1[2355], bank0[2355]} = 32'h0;
    {bank3[2356], bank2[2356], bank1[2356], bank0[2356]} = 32'h0;
    {bank3[2357], bank2[2357], bank1[2357], bank0[2357]} = 32'h0;
    {bank3[2358], bank2[2358], bank1[2358], bank0[2358]} = 32'h0;
    {bank3[2359], bank2[2359], bank1[2359], bank0[2359]} = 32'h0;
    {bank3[2360], bank2[2360], bank1[2360], bank0[2360]} = 32'h0;
    {bank3[2361], bank2[2361], bank1[2361], bank0[2361]} = 32'h0;
    {bank3[2362], bank2[2362], bank1[2362], bank0[2362]} = 32'h0;
    {bank3[2363], bank2[2363], bank1[2363], bank0[2363]} = 32'h0;
    {bank3[2364], bank2[2364], bank1[2364], bank0[2364]} = 32'h0;
    {bank3[2365], bank2[2365], bank1[2365], bank0[2365]} = 32'h0;
    {bank3[2366], bank2[2366], bank1[2366], bank0[2366]} = 32'h0;
    {bank3[2367], bank2[2367], bank1[2367], bank0[2367]} = 32'h0;
    {bank3[2368], bank2[2368], bank1[2368], bank0[2368]} = 32'h0;
    {bank3[2369], bank2[2369], bank1[2369], bank0[2369]} = 32'h0;
    {bank3[2370], bank2[2370], bank1[2370], bank0[2370]} = 32'h0;
    {bank3[2371], bank2[2371], bank1[2371], bank0[2371]} = 32'h0;
    {bank3[2372], bank2[2372], bank1[2372], bank0[2372]} = 32'h0;
    {bank3[2373], bank2[2373], bank1[2373], bank0[2373]} = 32'h0;
    {bank3[2374], bank2[2374], bank1[2374], bank0[2374]} = 32'h0;
    {bank3[2375], bank2[2375], bank1[2375], bank0[2375]} = 32'h0;
    {bank3[2376], bank2[2376], bank1[2376], bank0[2376]} = 32'h0;
    {bank3[2377], bank2[2377], bank1[2377], bank0[2377]} = 32'h0;
    {bank3[2378], bank2[2378], bank1[2378], bank0[2378]} = 32'h0;
    {bank3[2379], bank2[2379], bank1[2379], bank0[2379]} = 32'h0;
    {bank3[2380], bank2[2380], bank1[2380], bank0[2380]} = 32'h0;
    {bank3[2381], bank2[2381], bank1[2381], bank0[2381]} = 32'h0;
    {bank3[2382], bank2[2382], bank1[2382], bank0[2382]} = 32'h0;
    {bank3[2383], bank2[2383], bank1[2383], bank0[2383]} = 32'h0;
    {bank3[2384], bank2[2384], bank1[2384], bank0[2384]} = 32'h0;
    {bank3[2385], bank2[2385], bank1[2385], bank0[2385]} = 32'h0;
    {bank3[2386], bank2[2386], bank1[2386], bank0[2386]} = 32'h0;
    {bank3[2387], bank2[2387], bank1[2387], bank0[2387]} = 32'h0;
    {bank3[2388], bank2[2388], bank1[2388], bank0[2388]} = 32'h0;
    {bank3[2389], bank2[2389], bank1[2389], bank0[2389]} = 32'h0;
    {bank3[2390], bank2[2390], bank1[2390], bank0[2390]} = 32'h0;
    {bank3[2391], bank2[2391], bank1[2391], bank0[2391]} = 32'h0;
    {bank3[2392], bank2[2392], bank1[2392], bank0[2392]} = 32'h0;
    {bank3[2393], bank2[2393], bank1[2393], bank0[2393]} = 32'h0;
    {bank3[2394], bank2[2394], bank1[2394], bank0[2394]} = 32'h0;
    {bank3[2395], bank2[2395], bank1[2395], bank0[2395]} = 32'h0;
    {bank3[2396], bank2[2396], bank1[2396], bank0[2396]} = 32'h0;
    {bank3[2397], bank2[2397], bank1[2397], bank0[2397]} = 32'h0;
    {bank3[2398], bank2[2398], bank1[2398], bank0[2398]} = 32'h0;
    {bank3[2399], bank2[2399], bank1[2399], bank0[2399]} = 32'h0;
    {bank3[2400], bank2[2400], bank1[2400], bank0[2400]} = 32'h0;
    {bank3[2401], bank2[2401], bank1[2401], bank0[2401]} = 32'h0;
    {bank3[2402], bank2[2402], bank1[2402], bank0[2402]} = 32'h0;
    {bank3[2403], bank2[2403], bank1[2403], bank0[2403]} = 32'h0;
    {bank3[2404], bank2[2404], bank1[2404], bank0[2404]} = 32'h0;
    {bank3[2405], bank2[2405], bank1[2405], bank0[2405]} = 32'h0;
    {bank3[2406], bank2[2406], bank1[2406], bank0[2406]} = 32'h0;
    {bank3[2407], bank2[2407], bank1[2407], bank0[2407]} = 32'h0;
    {bank3[2408], bank2[2408], bank1[2408], bank0[2408]} = 32'h0;
    {bank3[2409], bank2[2409], bank1[2409], bank0[2409]} = 32'h0;
    {bank3[2410], bank2[2410], bank1[2410], bank0[2410]} = 32'h0;
    {bank3[2411], bank2[2411], bank1[2411], bank0[2411]} = 32'h0;
    {bank3[2412], bank2[2412], bank1[2412], bank0[2412]} = 32'h0;
    {bank3[2413], bank2[2413], bank1[2413], bank0[2413]} = 32'h0;
    {bank3[2414], bank2[2414], bank1[2414], bank0[2414]} = 32'h0;
    {bank3[2415], bank2[2415], bank1[2415], bank0[2415]} = 32'h0;
    {bank3[2416], bank2[2416], bank1[2416], bank0[2416]} = 32'h0;
    {bank3[2417], bank2[2417], bank1[2417], bank0[2417]} = 32'h0;
    {bank3[2418], bank2[2418], bank1[2418], bank0[2418]} = 32'h0;
    {bank3[2419], bank2[2419], bank1[2419], bank0[2419]} = 32'h0;
    {bank3[2420], bank2[2420], bank1[2420], bank0[2420]} = 32'h0;
    {bank3[2421], bank2[2421], bank1[2421], bank0[2421]} = 32'h0;
    {bank3[2422], bank2[2422], bank1[2422], bank0[2422]} = 32'h0;
    {bank3[2423], bank2[2423], bank1[2423], bank0[2423]} = 32'h0;
    {bank3[2424], bank2[2424], bank1[2424], bank0[2424]} = 32'h0;
    {bank3[2425], bank2[2425], bank1[2425], bank0[2425]} = 32'h0;
    {bank3[2426], bank2[2426], bank1[2426], bank0[2426]} = 32'h0;
    {bank3[2427], bank2[2427], bank1[2427], bank0[2427]} = 32'h0;
    {bank3[2428], bank2[2428], bank1[2428], bank0[2428]} = 32'h0;
    {bank3[2429], bank2[2429], bank1[2429], bank0[2429]} = 32'h0;
    {bank3[2430], bank2[2430], bank1[2430], bank0[2430]} = 32'h0;
    {bank3[2431], bank2[2431], bank1[2431], bank0[2431]} = 32'h0;
    {bank3[2432], bank2[2432], bank1[2432], bank0[2432]} = 32'h0;
    {bank3[2433], bank2[2433], bank1[2433], bank0[2433]} = 32'h0;
    {bank3[2434], bank2[2434], bank1[2434], bank0[2434]} = 32'h0;
    {bank3[2435], bank2[2435], bank1[2435], bank0[2435]} = 32'h0;
    {bank3[2436], bank2[2436], bank1[2436], bank0[2436]} = 32'h0;
    {bank3[2437], bank2[2437], bank1[2437], bank0[2437]} = 32'h0;
    {bank3[2438], bank2[2438], bank1[2438], bank0[2438]} = 32'h0;
    {bank3[2439], bank2[2439], bank1[2439], bank0[2439]} = 32'h0;
    {bank3[2440], bank2[2440], bank1[2440], bank0[2440]} = 32'h0;
    {bank3[2441], bank2[2441], bank1[2441], bank0[2441]} = 32'h0;
    {bank3[2442], bank2[2442], bank1[2442], bank0[2442]} = 32'h0;
    {bank3[2443], bank2[2443], bank1[2443], bank0[2443]} = 32'h0;
    {bank3[2444], bank2[2444], bank1[2444], bank0[2444]} = 32'h0;
    {bank3[2445], bank2[2445], bank1[2445], bank0[2445]} = 32'h0;
    {bank3[2446], bank2[2446], bank1[2446], bank0[2446]} = 32'h0;
    {bank3[2447], bank2[2447], bank1[2447], bank0[2447]} = 32'h0;
    {bank3[2448], bank2[2448], bank1[2448], bank0[2448]} = 32'h0;
    {bank3[2449], bank2[2449], bank1[2449], bank0[2449]} = 32'h0;
    {bank3[2450], bank2[2450], bank1[2450], bank0[2450]} = 32'h0;
    {bank3[2451], bank2[2451], bank1[2451], bank0[2451]} = 32'h0;
    {bank3[2452], bank2[2452], bank1[2452], bank0[2452]} = 32'h0;
    {bank3[2453], bank2[2453], bank1[2453], bank0[2453]} = 32'h0;
    {bank3[2454], bank2[2454], bank1[2454], bank0[2454]} = 32'h0;
    {bank3[2455], bank2[2455], bank1[2455], bank0[2455]} = 32'h0;
    {bank3[2456], bank2[2456], bank1[2456], bank0[2456]} = 32'h0;
    {bank3[2457], bank2[2457], bank1[2457], bank0[2457]} = 32'h0;
    {bank3[2458], bank2[2458], bank1[2458], bank0[2458]} = 32'h0;
    {bank3[2459], bank2[2459], bank1[2459], bank0[2459]} = 32'h0;
    {bank3[2460], bank2[2460], bank1[2460], bank0[2460]} = 32'h0;
    {bank3[2461], bank2[2461], bank1[2461], bank0[2461]} = 32'h0;
    {bank3[2462], bank2[2462], bank1[2462], bank0[2462]} = 32'h0;
    {bank3[2463], bank2[2463], bank1[2463], bank0[2463]} = 32'h0;
    {bank3[2464], bank2[2464], bank1[2464], bank0[2464]} = 32'h0;
    {bank3[2465], bank2[2465], bank1[2465], bank0[2465]} = 32'h0;
    {bank3[2466], bank2[2466], bank1[2466], bank0[2466]} = 32'h0;
    {bank3[2467], bank2[2467], bank1[2467], bank0[2467]} = 32'h0;
    {bank3[2468], bank2[2468], bank1[2468], bank0[2468]} = 32'h0;
    {bank3[2469], bank2[2469], bank1[2469], bank0[2469]} = 32'h0;
    {bank3[2470], bank2[2470], bank1[2470], bank0[2470]} = 32'h0;
    {bank3[2471], bank2[2471], bank1[2471], bank0[2471]} = 32'h0;
    {bank3[2472], bank2[2472], bank1[2472], bank0[2472]} = 32'h0;
    {bank3[2473], bank2[2473], bank1[2473], bank0[2473]} = 32'h0;
    {bank3[2474], bank2[2474], bank1[2474], bank0[2474]} = 32'h0;
    {bank3[2475], bank2[2475], bank1[2475], bank0[2475]} = 32'h0;
    {bank3[2476], bank2[2476], bank1[2476], bank0[2476]} = 32'h0;
    {bank3[2477], bank2[2477], bank1[2477], bank0[2477]} = 32'h0;
    {bank3[2478], bank2[2478], bank1[2478], bank0[2478]} = 32'h0;
    {bank3[2479], bank2[2479], bank1[2479], bank0[2479]} = 32'h0;
    {bank3[2480], bank2[2480], bank1[2480], bank0[2480]} = 32'h0;
    {bank3[2481], bank2[2481], bank1[2481], bank0[2481]} = 32'h0;
    {bank3[2482], bank2[2482], bank1[2482], bank0[2482]} = 32'h0;
    {bank3[2483], bank2[2483], bank1[2483], bank0[2483]} = 32'h0;
    {bank3[2484], bank2[2484], bank1[2484], bank0[2484]} = 32'h0;
    {bank3[2485], bank2[2485], bank1[2485], bank0[2485]} = 32'h0;
    {bank3[2486], bank2[2486], bank1[2486], bank0[2486]} = 32'h0;
    {bank3[2487], bank2[2487], bank1[2487], bank0[2487]} = 32'h0;
    {bank3[2488], bank2[2488], bank1[2488], bank0[2488]} = 32'h0;
    {bank3[2489], bank2[2489], bank1[2489], bank0[2489]} = 32'h0;
    {bank3[2490], bank2[2490], bank1[2490], bank0[2490]} = 32'h0;
    {bank3[2491], bank2[2491], bank1[2491], bank0[2491]} = 32'h0;
    {bank3[2492], bank2[2492], bank1[2492], bank0[2492]} = 32'h0;
    {bank3[2493], bank2[2493], bank1[2493], bank0[2493]} = 32'h0;
    {bank3[2494], bank2[2494], bank1[2494], bank0[2494]} = 32'h0;
    {bank3[2495], bank2[2495], bank1[2495], bank0[2495]} = 32'h0;
    {bank3[2496], bank2[2496], bank1[2496], bank0[2496]} = 32'h0;
    {bank3[2497], bank2[2497], bank1[2497], bank0[2497]} = 32'h0;
    {bank3[2498], bank2[2498], bank1[2498], bank0[2498]} = 32'h0;
    {bank3[2499], bank2[2499], bank1[2499], bank0[2499]} = 32'h0;
    {bank3[2500], bank2[2500], bank1[2500], bank0[2500]} = 32'h0;
    {bank3[2501], bank2[2501], bank1[2501], bank0[2501]} = 32'h0;
    {bank3[2502], bank2[2502], bank1[2502], bank0[2502]} = 32'h0;
    {bank3[2503], bank2[2503], bank1[2503], bank0[2503]} = 32'h0;
    {bank3[2504], bank2[2504], bank1[2504], bank0[2504]} = 32'h0;
    {bank3[2505], bank2[2505], bank1[2505], bank0[2505]} = 32'h0;
    {bank3[2506], bank2[2506], bank1[2506], bank0[2506]} = 32'h0;
    {bank3[2507], bank2[2507], bank1[2507], bank0[2507]} = 32'h0;
    {bank3[2508], bank2[2508], bank1[2508], bank0[2508]} = 32'h0;
    {bank3[2509], bank2[2509], bank1[2509], bank0[2509]} = 32'h0;
    {bank3[2510], bank2[2510], bank1[2510], bank0[2510]} = 32'h0;
    {bank3[2511], bank2[2511], bank1[2511], bank0[2511]} = 32'h0;
    {bank3[2512], bank2[2512], bank1[2512], bank0[2512]} = 32'h0;
    {bank3[2513], bank2[2513], bank1[2513], bank0[2513]} = 32'h0;
    {bank3[2514], bank2[2514], bank1[2514], bank0[2514]} = 32'h0;
    {bank3[2515], bank2[2515], bank1[2515], bank0[2515]} = 32'h0;
    {bank3[2516], bank2[2516], bank1[2516], bank0[2516]} = 32'h0;
    {bank3[2517], bank2[2517], bank1[2517], bank0[2517]} = 32'h0;
    {bank3[2518], bank2[2518], bank1[2518], bank0[2518]} = 32'h0;
    {bank3[2519], bank2[2519], bank1[2519], bank0[2519]} = 32'h0;
    {bank3[2520], bank2[2520], bank1[2520], bank0[2520]} = 32'h0;
    {bank3[2521], bank2[2521], bank1[2521], bank0[2521]} = 32'h0;
    {bank3[2522], bank2[2522], bank1[2522], bank0[2522]} = 32'h0;
    {bank3[2523], bank2[2523], bank1[2523], bank0[2523]} = 32'h0;
    {bank3[2524], bank2[2524], bank1[2524], bank0[2524]} = 32'h0;
    {bank3[2525], bank2[2525], bank1[2525], bank0[2525]} = 32'h0;
    {bank3[2526], bank2[2526], bank1[2526], bank0[2526]} = 32'h0;
    {bank3[2527], bank2[2527], bank1[2527], bank0[2527]} = 32'h0;
    {bank3[2528], bank2[2528], bank1[2528], bank0[2528]} = 32'h0;
    {bank3[2529], bank2[2529], bank1[2529], bank0[2529]} = 32'h0;
    {bank3[2530], bank2[2530], bank1[2530], bank0[2530]} = 32'h0;
    {bank3[2531], bank2[2531], bank1[2531], bank0[2531]} = 32'h0;
    {bank3[2532], bank2[2532], bank1[2532], bank0[2532]} = 32'h0;
    {bank3[2533], bank2[2533], bank1[2533], bank0[2533]} = 32'h0;
    {bank3[2534], bank2[2534], bank1[2534], bank0[2534]} = 32'h0;
    {bank3[2535], bank2[2535], bank1[2535], bank0[2535]} = 32'h0;
    {bank3[2536], bank2[2536], bank1[2536], bank0[2536]} = 32'h0;
    {bank3[2537], bank2[2537], bank1[2537], bank0[2537]} = 32'h0;
    {bank3[2538], bank2[2538], bank1[2538], bank0[2538]} = 32'h0;
    {bank3[2539], bank2[2539], bank1[2539], bank0[2539]} = 32'h0;
    {bank3[2540], bank2[2540], bank1[2540], bank0[2540]} = 32'h0;
    {bank3[2541], bank2[2541], bank1[2541], bank0[2541]} = 32'h0;
    {bank3[2542], bank2[2542], bank1[2542], bank0[2542]} = 32'h0;
    {bank3[2543], bank2[2543], bank1[2543], bank0[2543]} = 32'h0;
    {bank3[2544], bank2[2544], bank1[2544], bank0[2544]} = 32'h0;
    {bank3[2545], bank2[2545], bank1[2545], bank0[2545]} = 32'h0;
    {bank3[2546], bank2[2546], bank1[2546], bank0[2546]} = 32'h0;
    {bank3[2547], bank2[2547], bank1[2547], bank0[2547]} = 32'h0;
    {bank3[2548], bank2[2548], bank1[2548], bank0[2548]} = 32'h0;
    {bank3[2549], bank2[2549], bank1[2549], bank0[2549]} = 32'h0;
    {bank3[2550], bank2[2550], bank1[2550], bank0[2550]} = 32'h0;
    {bank3[2551], bank2[2551], bank1[2551], bank0[2551]} = 32'h0;
    {bank3[2552], bank2[2552], bank1[2552], bank0[2552]} = 32'h0;
    {bank3[2553], bank2[2553], bank1[2553], bank0[2553]} = 32'h0;
    {bank3[2554], bank2[2554], bank1[2554], bank0[2554]} = 32'h0;
    {bank3[2555], bank2[2555], bank1[2555], bank0[2555]} = 32'h0;
    {bank3[2556], bank2[2556], bank1[2556], bank0[2556]} = 32'h0;
    {bank3[2557], bank2[2557], bank1[2557], bank0[2557]} = 32'h0;
    {bank3[2558], bank2[2558], bank1[2558], bank0[2558]} = 32'h0;
    {bank3[2559], bank2[2559], bank1[2559], bank0[2559]} = 32'h0;
    {bank3[2560], bank2[2560], bank1[2560], bank0[2560]} = 32'h0;
    {bank3[2561], bank2[2561], bank1[2561], bank0[2561]} = 32'h0;
    {bank3[2562], bank2[2562], bank1[2562], bank0[2562]} = 32'h0;
    {bank3[2563], bank2[2563], bank1[2563], bank0[2563]} = 32'h0;
    {bank3[2564], bank2[2564], bank1[2564], bank0[2564]} = 32'h0;
    {bank3[2565], bank2[2565], bank1[2565], bank0[2565]} = 32'h0;
    {bank3[2566], bank2[2566], bank1[2566], bank0[2566]} = 32'h0;
    {bank3[2567], bank2[2567], bank1[2567], bank0[2567]} = 32'h0;
    {bank3[2568], bank2[2568], bank1[2568], bank0[2568]} = 32'h0;
    {bank3[2569], bank2[2569], bank1[2569], bank0[2569]} = 32'h0;
    {bank3[2570], bank2[2570], bank1[2570], bank0[2570]} = 32'h0;
    {bank3[2571], bank2[2571], bank1[2571], bank0[2571]} = 32'h0;
    {bank3[2572], bank2[2572], bank1[2572], bank0[2572]} = 32'h0;
    {bank3[2573], bank2[2573], bank1[2573], bank0[2573]} = 32'h0;
    {bank3[2574], bank2[2574], bank1[2574], bank0[2574]} = 32'h0;
    {bank3[2575], bank2[2575], bank1[2575], bank0[2575]} = 32'h0;
    {bank3[2576], bank2[2576], bank1[2576], bank0[2576]} = 32'h0;
    {bank3[2577], bank2[2577], bank1[2577], bank0[2577]} = 32'h0;
    {bank3[2578], bank2[2578], bank1[2578], bank0[2578]} = 32'h0;
    {bank3[2579], bank2[2579], bank1[2579], bank0[2579]} = 32'h0;
    {bank3[2580], bank2[2580], bank1[2580], bank0[2580]} = 32'h0;
    {bank3[2581], bank2[2581], bank1[2581], bank0[2581]} = 32'h0;
    {bank3[2582], bank2[2582], bank1[2582], bank0[2582]} = 32'h0;
    {bank3[2583], bank2[2583], bank1[2583], bank0[2583]} = 32'h0;
    {bank3[2584], bank2[2584], bank1[2584], bank0[2584]} = 32'h0;
    {bank3[2585], bank2[2585], bank1[2585], bank0[2585]} = 32'h0;
    {bank3[2586], bank2[2586], bank1[2586], bank0[2586]} = 32'h0;
    {bank3[2587], bank2[2587], bank1[2587], bank0[2587]} = 32'h0;
    {bank3[2588], bank2[2588], bank1[2588], bank0[2588]} = 32'h0;
    {bank3[2589], bank2[2589], bank1[2589], bank0[2589]} = 32'h0;
    {bank3[2590], bank2[2590], bank1[2590], bank0[2590]} = 32'h0;
    {bank3[2591], bank2[2591], bank1[2591], bank0[2591]} = 32'h0;
    {bank3[2592], bank2[2592], bank1[2592], bank0[2592]} = 32'h0;
    {bank3[2593], bank2[2593], bank1[2593], bank0[2593]} = 32'h0;
    {bank3[2594], bank2[2594], bank1[2594], bank0[2594]} = 32'h0;
    {bank3[2595], bank2[2595], bank1[2595], bank0[2595]} = 32'h0;
    {bank3[2596], bank2[2596], bank1[2596], bank0[2596]} = 32'h0;
    {bank3[2597], bank2[2597], bank1[2597], bank0[2597]} = 32'h0;
    {bank3[2598], bank2[2598], bank1[2598], bank0[2598]} = 32'h0;
    {bank3[2599], bank2[2599], bank1[2599], bank0[2599]} = 32'h0;
    {bank3[2600], bank2[2600], bank1[2600], bank0[2600]} = 32'h0;
    {bank3[2601], bank2[2601], bank1[2601], bank0[2601]} = 32'h0;
    {bank3[2602], bank2[2602], bank1[2602], bank0[2602]} = 32'h0;
    {bank3[2603], bank2[2603], bank1[2603], bank0[2603]} = 32'h0;
    {bank3[2604], bank2[2604], bank1[2604], bank0[2604]} = 32'h0;
    {bank3[2605], bank2[2605], bank1[2605], bank0[2605]} = 32'h0;
    {bank3[2606], bank2[2606], bank1[2606], bank0[2606]} = 32'h0;
    {bank3[2607], bank2[2607], bank1[2607], bank0[2607]} = 32'h0;
    {bank3[2608], bank2[2608], bank1[2608], bank0[2608]} = 32'h0;
    {bank3[2609], bank2[2609], bank1[2609], bank0[2609]} = 32'h0;
    {bank3[2610], bank2[2610], bank1[2610], bank0[2610]} = 32'h0;
    {bank3[2611], bank2[2611], bank1[2611], bank0[2611]} = 32'h0;
    {bank3[2612], bank2[2612], bank1[2612], bank0[2612]} = 32'h0;
    {bank3[2613], bank2[2613], bank1[2613], bank0[2613]} = 32'h0;
    {bank3[2614], bank2[2614], bank1[2614], bank0[2614]} = 32'h0;
    {bank3[2615], bank2[2615], bank1[2615], bank0[2615]} = 32'h0;
    {bank3[2616], bank2[2616], bank1[2616], bank0[2616]} = 32'h0;
    {bank3[2617], bank2[2617], bank1[2617], bank0[2617]} = 32'h0;
    {bank3[2618], bank2[2618], bank1[2618], bank0[2618]} = 32'h0;
    {bank3[2619], bank2[2619], bank1[2619], bank0[2619]} = 32'h0;
    {bank3[2620], bank2[2620], bank1[2620], bank0[2620]} = 32'h0;
    {bank3[2621], bank2[2621], bank1[2621], bank0[2621]} = 32'h0;
    {bank3[2622], bank2[2622], bank1[2622], bank0[2622]} = 32'h0;
    {bank3[2623], bank2[2623], bank1[2623], bank0[2623]} = 32'h0;
    {bank3[2624], bank2[2624], bank1[2624], bank0[2624]} = 32'h0;
    {bank3[2625], bank2[2625], bank1[2625], bank0[2625]} = 32'h0;
    {bank3[2626], bank2[2626], bank1[2626], bank0[2626]} = 32'h0;
    {bank3[2627], bank2[2627], bank1[2627], bank0[2627]} = 32'h0;
    {bank3[2628], bank2[2628], bank1[2628], bank0[2628]} = 32'h0;
    {bank3[2629], bank2[2629], bank1[2629], bank0[2629]} = 32'h0;
    {bank3[2630], bank2[2630], bank1[2630], bank0[2630]} = 32'h0;
    {bank3[2631], bank2[2631], bank1[2631], bank0[2631]} = 32'h0;
    {bank3[2632], bank2[2632], bank1[2632], bank0[2632]} = 32'h0;
    {bank3[2633], bank2[2633], bank1[2633], bank0[2633]} = 32'h0;
    {bank3[2634], bank2[2634], bank1[2634], bank0[2634]} = 32'h0;
    {bank3[2635], bank2[2635], bank1[2635], bank0[2635]} = 32'h0;
    {bank3[2636], bank2[2636], bank1[2636], bank0[2636]} = 32'h0;
    {bank3[2637], bank2[2637], bank1[2637], bank0[2637]} = 32'h0;
    {bank3[2638], bank2[2638], bank1[2638], bank0[2638]} = 32'h0;
    {bank3[2639], bank2[2639], bank1[2639], bank0[2639]} = 32'h0;
    {bank3[2640], bank2[2640], bank1[2640], bank0[2640]} = 32'h0;
    {bank3[2641], bank2[2641], bank1[2641], bank0[2641]} = 32'h0;
    {bank3[2642], bank2[2642], bank1[2642], bank0[2642]} = 32'h0;
    {bank3[2643], bank2[2643], bank1[2643], bank0[2643]} = 32'h0;
    {bank3[2644], bank2[2644], bank1[2644], bank0[2644]} = 32'h0;
    {bank3[2645], bank2[2645], bank1[2645], bank0[2645]} = 32'h0;
    {bank3[2646], bank2[2646], bank1[2646], bank0[2646]} = 32'h0;
    {bank3[2647], bank2[2647], bank1[2647], bank0[2647]} = 32'h0;
    {bank3[2648], bank2[2648], bank1[2648], bank0[2648]} = 32'h0;
    {bank3[2649], bank2[2649], bank1[2649], bank0[2649]} = 32'h0;
    {bank3[2650], bank2[2650], bank1[2650], bank0[2650]} = 32'h0;
    {bank3[2651], bank2[2651], bank1[2651], bank0[2651]} = 32'h0;
    {bank3[2652], bank2[2652], bank1[2652], bank0[2652]} = 32'h0;
    {bank3[2653], bank2[2653], bank1[2653], bank0[2653]} = 32'h0;
    {bank3[2654], bank2[2654], bank1[2654], bank0[2654]} = 32'h0;
    {bank3[2655], bank2[2655], bank1[2655], bank0[2655]} = 32'h0;
    {bank3[2656], bank2[2656], bank1[2656], bank0[2656]} = 32'h0;
    {bank3[2657], bank2[2657], bank1[2657], bank0[2657]} = 32'h0;
    {bank3[2658], bank2[2658], bank1[2658], bank0[2658]} = 32'h0;
    {bank3[2659], bank2[2659], bank1[2659], bank0[2659]} = 32'h0;
    {bank3[2660], bank2[2660], bank1[2660], bank0[2660]} = 32'h0;
    {bank3[2661], bank2[2661], bank1[2661], bank0[2661]} = 32'h0;
    {bank3[2662], bank2[2662], bank1[2662], bank0[2662]} = 32'h0;
    {bank3[2663], bank2[2663], bank1[2663], bank0[2663]} = 32'h0;
    {bank3[2664], bank2[2664], bank1[2664], bank0[2664]} = 32'h0;
    {bank3[2665], bank2[2665], bank1[2665], bank0[2665]} = 32'h0;
    {bank3[2666], bank2[2666], bank1[2666], bank0[2666]} = 32'h0;
    {bank3[2667], bank2[2667], bank1[2667], bank0[2667]} = 32'h0;
    {bank3[2668], bank2[2668], bank1[2668], bank0[2668]} = 32'h0;
    {bank3[2669], bank2[2669], bank1[2669], bank0[2669]} = 32'h0;
    {bank3[2670], bank2[2670], bank1[2670], bank0[2670]} = 32'h0;
    {bank3[2671], bank2[2671], bank1[2671], bank0[2671]} = 32'h0;
    {bank3[2672], bank2[2672], bank1[2672], bank0[2672]} = 32'h0;
    {bank3[2673], bank2[2673], bank1[2673], bank0[2673]} = 32'h0;
    {bank3[2674], bank2[2674], bank1[2674], bank0[2674]} = 32'h0;
    {bank3[2675], bank2[2675], bank1[2675], bank0[2675]} = 32'h0;
    {bank3[2676], bank2[2676], bank1[2676], bank0[2676]} = 32'h0;
    {bank3[2677], bank2[2677], bank1[2677], bank0[2677]} = 32'h0;
    {bank3[2678], bank2[2678], bank1[2678], bank0[2678]} = 32'h0;
    {bank3[2679], bank2[2679], bank1[2679], bank0[2679]} = 32'h0;
    {bank3[2680], bank2[2680], bank1[2680], bank0[2680]} = 32'h0;
    {bank3[2681], bank2[2681], bank1[2681], bank0[2681]} = 32'h0;
    {bank3[2682], bank2[2682], bank1[2682], bank0[2682]} = 32'h0;
    {bank3[2683], bank2[2683], bank1[2683], bank0[2683]} = 32'h0;
    {bank3[2684], bank2[2684], bank1[2684], bank0[2684]} = 32'h0;
    {bank3[2685], bank2[2685], bank1[2685], bank0[2685]} = 32'h0;
    {bank3[2686], bank2[2686], bank1[2686], bank0[2686]} = 32'h0;
    {bank3[2687], bank2[2687], bank1[2687], bank0[2687]} = 32'h0;
    {bank3[2688], bank2[2688], bank1[2688], bank0[2688]} = 32'h0;
    {bank3[2689], bank2[2689], bank1[2689], bank0[2689]} = 32'h0;
    {bank3[2690], bank2[2690], bank1[2690], bank0[2690]} = 32'h0;
    {bank3[2691], bank2[2691], bank1[2691], bank0[2691]} = 32'h0;
    {bank3[2692], bank2[2692], bank1[2692], bank0[2692]} = 32'h0;
    {bank3[2693], bank2[2693], bank1[2693], bank0[2693]} = 32'h0;
    {bank3[2694], bank2[2694], bank1[2694], bank0[2694]} = 32'h0;
    {bank3[2695], bank2[2695], bank1[2695], bank0[2695]} = 32'h0;
    {bank3[2696], bank2[2696], bank1[2696], bank0[2696]} = 32'h0;
    {bank3[2697], bank2[2697], bank1[2697], bank0[2697]} = 32'h0;
    {bank3[2698], bank2[2698], bank1[2698], bank0[2698]} = 32'h0;
    {bank3[2699], bank2[2699], bank1[2699], bank0[2699]} = 32'h0;
    {bank3[2700], bank2[2700], bank1[2700], bank0[2700]} = 32'h0;
    {bank3[2701], bank2[2701], bank1[2701], bank0[2701]} = 32'h0;
    {bank3[2702], bank2[2702], bank1[2702], bank0[2702]} = 32'h0;
    {bank3[2703], bank2[2703], bank1[2703], bank0[2703]} = 32'h0;
    {bank3[2704], bank2[2704], bank1[2704], bank0[2704]} = 32'h0;
    {bank3[2705], bank2[2705], bank1[2705], bank0[2705]} = 32'h0;
    {bank3[2706], bank2[2706], bank1[2706], bank0[2706]} = 32'h0;
    {bank3[2707], bank2[2707], bank1[2707], bank0[2707]} = 32'h0;
    {bank3[2708], bank2[2708], bank1[2708], bank0[2708]} = 32'h0;
    {bank3[2709], bank2[2709], bank1[2709], bank0[2709]} = 32'h0;
    {bank3[2710], bank2[2710], bank1[2710], bank0[2710]} = 32'h0;
    {bank3[2711], bank2[2711], bank1[2711], bank0[2711]} = 32'h0;
    {bank3[2712], bank2[2712], bank1[2712], bank0[2712]} = 32'h0;
    {bank3[2713], bank2[2713], bank1[2713], bank0[2713]} = 32'h0;
    {bank3[2714], bank2[2714], bank1[2714], bank0[2714]} = 32'h0;
    {bank3[2715], bank2[2715], bank1[2715], bank0[2715]} = 32'h0;
    {bank3[2716], bank2[2716], bank1[2716], bank0[2716]} = 32'h0;
    {bank3[2717], bank2[2717], bank1[2717], bank0[2717]} = 32'h0;
    {bank3[2718], bank2[2718], bank1[2718], bank0[2718]} = 32'h0;
    {bank3[2719], bank2[2719], bank1[2719], bank0[2719]} = 32'h0;
    {bank3[2720], bank2[2720], bank1[2720], bank0[2720]} = 32'h0;
    {bank3[2721], bank2[2721], bank1[2721], bank0[2721]} = 32'h0;
    {bank3[2722], bank2[2722], bank1[2722], bank0[2722]} = 32'h0;
    {bank3[2723], bank2[2723], bank1[2723], bank0[2723]} = 32'h0;
    {bank3[2724], bank2[2724], bank1[2724], bank0[2724]} = 32'h0;
    {bank3[2725], bank2[2725], bank1[2725], bank0[2725]} = 32'h0;
    {bank3[2726], bank2[2726], bank1[2726], bank0[2726]} = 32'h0;
    {bank3[2727], bank2[2727], bank1[2727], bank0[2727]} = 32'h0;
    {bank3[2728], bank2[2728], bank1[2728], bank0[2728]} = 32'h0;
    {bank3[2729], bank2[2729], bank1[2729], bank0[2729]} = 32'h0;
    {bank3[2730], bank2[2730], bank1[2730], bank0[2730]} = 32'h0;
    {bank3[2731], bank2[2731], bank1[2731], bank0[2731]} = 32'h0;
    {bank3[2732], bank2[2732], bank1[2732], bank0[2732]} = 32'h0;
    {bank3[2733], bank2[2733], bank1[2733], bank0[2733]} = 32'h0;
    {bank3[2734], bank2[2734], bank1[2734], bank0[2734]} = 32'h0;
    {bank3[2735], bank2[2735], bank1[2735], bank0[2735]} = 32'h0;
    {bank3[2736], bank2[2736], bank1[2736], bank0[2736]} = 32'h0;
    {bank3[2737], bank2[2737], bank1[2737], bank0[2737]} = 32'h0;
    {bank3[2738], bank2[2738], bank1[2738], bank0[2738]} = 32'h0;
    {bank3[2739], bank2[2739], bank1[2739], bank0[2739]} = 32'h0;
    {bank3[2740], bank2[2740], bank1[2740], bank0[2740]} = 32'h0;
    {bank3[2741], bank2[2741], bank1[2741], bank0[2741]} = 32'h0;
    {bank3[2742], bank2[2742], bank1[2742], bank0[2742]} = 32'h0;
    {bank3[2743], bank2[2743], bank1[2743], bank0[2743]} = 32'h0;
    {bank3[2744], bank2[2744], bank1[2744], bank0[2744]} = 32'h0;
    {bank3[2745], bank2[2745], bank1[2745], bank0[2745]} = 32'h0;
    {bank3[2746], bank2[2746], bank1[2746], bank0[2746]} = 32'h0;
    {bank3[2747], bank2[2747], bank1[2747], bank0[2747]} = 32'h0;
    {bank3[2748], bank2[2748], bank1[2748], bank0[2748]} = 32'h0;
    {bank3[2749], bank2[2749], bank1[2749], bank0[2749]} = 32'h0;
    {bank3[2750], bank2[2750], bank1[2750], bank0[2750]} = 32'h0;
    {bank3[2751], bank2[2751], bank1[2751], bank0[2751]} = 32'h0;
    {bank3[2752], bank2[2752], bank1[2752], bank0[2752]} = 32'h0;
    {bank3[2753], bank2[2753], bank1[2753], bank0[2753]} = 32'h0;
    {bank3[2754], bank2[2754], bank1[2754], bank0[2754]} = 32'h0;
    {bank3[2755], bank2[2755], bank1[2755], bank0[2755]} = 32'h0;
    {bank3[2756], bank2[2756], bank1[2756], bank0[2756]} = 32'h0;
    {bank3[2757], bank2[2757], bank1[2757], bank0[2757]} = 32'h0;
    {bank3[2758], bank2[2758], bank1[2758], bank0[2758]} = 32'h0;
    {bank3[2759], bank2[2759], bank1[2759], bank0[2759]} = 32'h0;
    {bank3[2760], bank2[2760], bank1[2760], bank0[2760]} = 32'h0;
    {bank3[2761], bank2[2761], bank1[2761], bank0[2761]} = 32'h0;
    {bank3[2762], bank2[2762], bank1[2762], bank0[2762]} = 32'h0;
    {bank3[2763], bank2[2763], bank1[2763], bank0[2763]} = 32'h0;
    {bank3[2764], bank2[2764], bank1[2764], bank0[2764]} = 32'h0;
    {bank3[2765], bank2[2765], bank1[2765], bank0[2765]} = 32'h0;
    {bank3[2766], bank2[2766], bank1[2766], bank0[2766]} = 32'h0;
    {bank3[2767], bank2[2767], bank1[2767], bank0[2767]} = 32'h0;
    {bank3[2768], bank2[2768], bank1[2768], bank0[2768]} = 32'h0;
    {bank3[2769], bank2[2769], bank1[2769], bank0[2769]} = 32'h0;
    {bank3[2770], bank2[2770], bank1[2770], bank0[2770]} = 32'h0;
    {bank3[2771], bank2[2771], bank1[2771], bank0[2771]} = 32'h0;
    {bank3[2772], bank2[2772], bank1[2772], bank0[2772]} = 32'h0;
    {bank3[2773], bank2[2773], bank1[2773], bank0[2773]} = 32'h0;
    {bank3[2774], bank2[2774], bank1[2774], bank0[2774]} = 32'h0;
    {bank3[2775], bank2[2775], bank1[2775], bank0[2775]} = 32'h0;
    {bank3[2776], bank2[2776], bank1[2776], bank0[2776]} = 32'h0;
    {bank3[2777], bank2[2777], bank1[2777], bank0[2777]} = 32'h0;
    {bank3[2778], bank2[2778], bank1[2778], bank0[2778]} = 32'h0;
    {bank3[2779], bank2[2779], bank1[2779], bank0[2779]} = 32'h0;
    {bank3[2780], bank2[2780], bank1[2780], bank0[2780]} = 32'h0;
    {bank3[2781], bank2[2781], bank1[2781], bank0[2781]} = 32'h0;
    {bank3[2782], bank2[2782], bank1[2782], bank0[2782]} = 32'h0;
    {bank3[2783], bank2[2783], bank1[2783], bank0[2783]} = 32'h0;
    {bank3[2784], bank2[2784], bank1[2784], bank0[2784]} = 32'h0;
    {bank3[2785], bank2[2785], bank1[2785], bank0[2785]} = 32'h0;
    {bank3[2786], bank2[2786], bank1[2786], bank0[2786]} = 32'h0;
    {bank3[2787], bank2[2787], bank1[2787], bank0[2787]} = 32'h0;
    {bank3[2788], bank2[2788], bank1[2788], bank0[2788]} = 32'h0;
    {bank3[2789], bank2[2789], bank1[2789], bank0[2789]} = 32'h0;
    {bank3[2790], bank2[2790], bank1[2790], bank0[2790]} = 32'h0;
    {bank3[2791], bank2[2791], bank1[2791], bank0[2791]} = 32'h0;
    {bank3[2792], bank2[2792], bank1[2792], bank0[2792]} = 32'h0;
    {bank3[2793], bank2[2793], bank1[2793], bank0[2793]} = 32'h0;
    {bank3[2794], bank2[2794], bank1[2794], bank0[2794]} = 32'h0;
    {bank3[2795], bank2[2795], bank1[2795], bank0[2795]} = 32'h0;
    {bank3[2796], bank2[2796], bank1[2796], bank0[2796]} = 32'h0;
    {bank3[2797], bank2[2797], bank1[2797], bank0[2797]} = 32'h0;
    {bank3[2798], bank2[2798], bank1[2798], bank0[2798]} = 32'h0;
    {bank3[2799], bank2[2799], bank1[2799], bank0[2799]} = 32'h0;
    {bank3[2800], bank2[2800], bank1[2800], bank0[2800]} = 32'h0;
    {bank3[2801], bank2[2801], bank1[2801], bank0[2801]} = 32'h0;
    {bank3[2802], bank2[2802], bank1[2802], bank0[2802]} = 32'h0;
    {bank3[2803], bank2[2803], bank1[2803], bank0[2803]} = 32'h0;
    {bank3[2804], bank2[2804], bank1[2804], bank0[2804]} = 32'h0;
    {bank3[2805], bank2[2805], bank1[2805], bank0[2805]} = 32'h0;
    {bank3[2806], bank2[2806], bank1[2806], bank0[2806]} = 32'h0;
    {bank3[2807], bank2[2807], bank1[2807], bank0[2807]} = 32'h0;
    {bank3[2808], bank2[2808], bank1[2808], bank0[2808]} = 32'h0;
    {bank3[2809], bank2[2809], bank1[2809], bank0[2809]} = 32'h0;
    {bank3[2810], bank2[2810], bank1[2810], bank0[2810]} = 32'h0;
    {bank3[2811], bank2[2811], bank1[2811], bank0[2811]} = 32'h0;
    {bank3[2812], bank2[2812], bank1[2812], bank0[2812]} = 32'h0;
    {bank3[2813], bank2[2813], bank1[2813], bank0[2813]} = 32'h0;
    {bank3[2814], bank2[2814], bank1[2814], bank0[2814]} = 32'h0;
    {bank3[2815], bank2[2815], bank1[2815], bank0[2815]} = 32'h0;
    {bank3[2816], bank2[2816], bank1[2816], bank0[2816]} = 32'h0;
    {bank3[2817], bank2[2817], bank1[2817], bank0[2817]} = 32'h0;
    {bank3[2818], bank2[2818], bank1[2818], bank0[2818]} = 32'h0;
    {bank3[2819], bank2[2819], bank1[2819], bank0[2819]} = 32'h0;
    {bank3[2820], bank2[2820], bank1[2820], bank0[2820]} = 32'h0;
    {bank3[2821], bank2[2821], bank1[2821], bank0[2821]} = 32'h0;
    {bank3[2822], bank2[2822], bank1[2822], bank0[2822]} = 32'h0;
    {bank3[2823], bank2[2823], bank1[2823], bank0[2823]} = 32'h0;
    {bank3[2824], bank2[2824], bank1[2824], bank0[2824]} = 32'h0;
    {bank3[2825], bank2[2825], bank1[2825], bank0[2825]} = 32'h0;
    {bank3[2826], bank2[2826], bank1[2826], bank0[2826]} = 32'h0;
    {bank3[2827], bank2[2827], bank1[2827], bank0[2827]} = 32'h0;
    {bank3[2828], bank2[2828], bank1[2828], bank0[2828]} = 32'h0;
    {bank3[2829], bank2[2829], bank1[2829], bank0[2829]} = 32'h0;
    {bank3[2830], bank2[2830], bank1[2830], bank0[2830]} = 32'h0;
    {bank3[2831], bank2[2831], bank1[2831], bank0[2831]} = 32'h0;
    {bank3[2832], bank2[2832], bank1[2832], bank0[2832]} = 32'h0;
    {bank3[2833], bank2[2833], bank1[2833], bank0[2833]} = 32'h0;
    {bank3[2834], bank2[2834], bank1[2834], bank0[2834]} = 32'h0;
    {bank3[2835], bank2[2835], bank1[2835], bank0[2835]} = 32'h0;
    {bank3[2836], bank2[2836], bank1[2836], bank0[2836]} = 32'h0;
    {bank3[2837], bank2[2837], bank1[2837], bank0[2837]} = 32'h0;
    {bank3[2838], bank2[2838], bank1[2838], bank0[2838]} = 32'h0;
    {bank3[2839], bank2[2839], bank1[2839], bank0[2839]} = 32'h0;
    {bank3[2840], bank2[2840], bank1[2840], bank0[2840]} = 32'h0;
    {bank3[2841], bank2[2841], bank1[2841], bank0[2841]} = 32'h0;
    {bank3[2842], bank2[2842], bank1[2842], bank0[2842]} = 32'h0;
    {bank3[2843], bank2[2843], bank1[2843], bank0[2843]} = 32'h0;
    {bank3[2844], bank2[2844], bank1[2844], bank0[2844]} = 32'h0;
    {bank3[2845], bank2[2845], bank1[2845], bank0[2845]} = 32'h0;
    {bank3[2846], bank2[2846], bank1[2846], bank0[2846]} = 32'h0;
    {bank3[2847], bank2[2847], bank1[2847], bank0[2847]} = 32'h0;
    {bank3[2848], bank2[2848], bank1[2848], bank0[2848]} = 32'h0;
    {bank3[2849], bank2[2849], bank1[2849], bank0[2849]} = 32'h0;
    {bank3[2850], bank2[2850], bank1[2850], bank0[2850]} = 32'h0;
    {bank3[2851], bank2[2851], bank1[2851], bank0[2851]} = 32'h0;
    {bank3[2852], bank2[2852], bank1[2852], bank0[2852]} = 32'h0;
    {bank3[2853], bank2[2853], bank1[2853], bank0[2853]} = 32'h0;
    {bank3[2854], bank2[2854], bank1[2854], bank0[2854]} = 32'h0;
    {bank3[2855], bank2[2855], bank1[2855], bank0[2855]} = 32'h0;
    {bank3[2856], bank2[2856], bank1[2856], bank0[2856]} = 32'h0;
    {bank3[2857], bank2[2857], bank1[2857], bank0[2857]} = 32'h0;
    {bank3[2858], bank2[2858], bank1[2858], bank0[2858]} = 32'h0;
    {bank3[2859], bank2[2859], bank1[2859], bank0[2859]} = 32'h0;
    {bank3[2860], bank2[2860], bank1[2860], bank0[2860]} = 32'h0;
    {bank3[2861], bank2[2861], bank1[2861], bank0[2861]} = 32'h0;
    {bank3[2862], bank2[2862], bank1[2862], bank0[2862]} = 32'h0;
    {bank3[2863], bank2[2863], bank1[2863], bank0[2863]} = 32'h0;
    {bank3[2864], bank2[2864], bank1[2864], bank0[2864]} = 32'h0;
    {bank3[2865], bank2[2865], bank1[2865], bank0[2865]} = 32'h0;
    {bank3[2866], bank2[2866], bank1[2866], bank0[2866]} = 32'h0;
    {bank3[2867], bank2[2867], bank1[2867], bank0[2867]} = 32'h0;
    {bank3[2868], bank2[2868], bank1[2868], bank0[2868]} = 32'h0;
    {bank3[2869], bank2[2869], bank1[2869], bank0[2869]} = 32'h0;
    {bank3[2870], bank2[2870], bank1[2870], bank0[2870]} = 32'h0;
    {bank3[2871], bank2[2871], bank1[2871], bank0[2871]} = 32'h0;
    {bank3[2872], bank2[2872], bank1[2872], bank0[2872]} = 32'h0;
    {bank3[2873], bank2[2873], bank1[2873], bank0[2873]} = 32'h0;
    {bank3[2874], bank2[2874], bank1[2874], bank0[2874]} = 32'h0;
    {bank3[2875], bank2[2875], bank1[2875], bank0[2875]} = 32'h0;
    {bank3[2876], bank2[2876], bank1[2876], bank0[2876]} = 32'h0;
    {bank3[2877], bank2[2877], bank1[2877], bank0[2877]} = 32'h0;
    {bank3[2878], bank2[2878], bank1[2878], bank0[2878]} = 32'h0;
    {bank3[2879], bank2[2879], bank1[2879], bank0[2879]} = 32'h0;
    {bank3[2880], bank2[2880], bank1[2880], bank0[2880]} = 32'h0;
    {bank3[2881], bank2[2881], bank1[2881], bank0[2881]} = 32'h0;
    {bank3[2882], bank2[2882], bank1[2882], bank0[2882]} = 32'h0;
    {bank3[2883], bank2[2883], bank1[2883], bank0[2883]} = 32'h0;
    {bank3[2884], bank2[2884], bank1[2884], bank0[2884]} = 32'h0;
    {bank3[2885], bank2[2885], bank1[2885], bank0[2885]} = 32'h0;
    {bank3[2886], bank2[2886], bank1[2886], bank0[2886]} = 32'h0;
    {bank3[2887], bank2[2887], bank1[2887], bank0[2887]} = 32'h0;
    {bank3[2888], bank2[2888], bank1[2888], bank0[2888]} = 32'h0;
    {bank3[2889], bank2[2889], bank1[2889], bank0[2889]} = 32'h0;
    {bank3[2890], bank2[2890], bank1[2890], bank0[2890]} = 32'h0;
    {bank3[2891], bank2[2891], bank1[2891], bank0[2891]} = 32'h0;
    {bank3[2892], bank2[2892], bank1[2892], bank0[2892]} = 32'h0;
    {bank3[2893], bank2[2893], bank1[2893], bank0[2893]} = 32'h0;
    {bank3[2894], bank2[2894], bank1[2894], bank0[2894]} = 32'h0;
    {bank3[2895], bank2[2895], bank1[2895], bank0[2895]} = 32'h0;
    {bank3[2896], bank2[2896], bank1[2896], bank0[2896]} = 32'h0;
    {bank3[2897], bank2[2897], bank1[2897], bank0[2897]} = 32'h0;
    {bank3[2898], bank2[2898], bank1[2898], bank0[2898]} = 32'h0;
    {bank3[2899], bank2[2899], bank1[2899], bank0[2899]} = 32'h0;
    {bank3[2900], bank2[2900], bank1[2900], bank0[2900]} = 32'h0;
    {bank3[2901], bank2[2901], bank1[2901], bank0[2901]} = 32'h0;
    {bank3[2902], bank2[2902], bank1[2902], bank0[2902]} = 32'h0;
    {bank3[2903], bank2[2903], bank1[2903], bank0[2903]} = 32'h0;
    {bank3[2904], bank2[2904], bank1[2904], bank0[2904]} = 32'h0;
    {bank3[2905], bank2[2905], bank1[2905], bank0[2905]} = 32'h0;
    {bank3[2906], bank2[2906], bank1[2906], bank0[2906]} = 32'h0;
    {bank3[2907], bank2[2907], bank1[2907], bank0[2907]} = 32'h0;
    {bank3[2908], bank2[2908], bank1[2908], bank0[2908]} = 32'h0;
    {bank3[2909], bank2[2909], bank1[2909], bank0[2909]} = 32'h0;
    {bank3[2910], bank2[2910], bank1[2910], bank0[2910]} = 32'h0;
    {bank3[2911], bank2[2911], bank1[2911], bank0[2911]} = 32'h0;
    {bank3[2912], bank2[2912], bank1[2912], bank0[2912]} = 32'h0;
    {bank3[2913], bank2[2913], bank1[2913], bank0[2913]} = 32'h0;
    {bank3[2914], bank2[2914], bank1[2914], bank0[2914]} = 32'h0;
    {bank3[2915], bank2[2915], bank1[2915], bank0[2915]} = 32'h0;
    {bank3[2916], bank2[2916], bank1[2916], bank0[2916]} = 32'h0;
    {bank3[2917], bank2[2917], bank1[2917], bank0[2917]} = 32'h0;
    {bank3[2918], bank2[2918], bank1[2918], bank0[2918]} = 32'h0;
    {bank3[2919], bank2[2919], bank1[2919], bank0[2919]} = 32'h0;
    {bank3[2920], bank2[2920], bank1[2920], bank0[2920]} = 32'h0;
    {bank3[2921], bank2[2921], bank1[2921], bank0[2921]} = 32'h0;
    {bank3[2922], bank2[2922], bank1[2922], bank0[2922]} = 32'h0;
    {bank3[2923], bank2[2923], bank1[2923], bank0[2923]} = 32'h0;
    {bank3[2924], bank2[2924], bank1[2924], bank0[2924]} = 32'h0;
    {bank3[2925], bank2[2925], bank1[2925], bank0[2925]} = 32'h0;
    {bank3[2926], bank2[2926], bank1[2926], bank0[2926]} = 32'h0;
    {bank3[2927], bank2[2927], bank1[2927], bank0[2927]} = 32'h0;
    {bank3[2928], bank2[2928], bank1[2928], bank0[2928]} = 32'h0;
    {bank3[2929], bank2[2929], bank1[2929], bank0[2929]} = 32'h0;
    {bank3[2930], bank2[2930], bank1[2930], bank0[2930]} = 32'h0;
    {bank3[2931], bank2[2931], bank1[2931], bank0[2931]} = 32'h0;
    {bank3[2932], bank2[2932], bank1[2932], bank0[2932]} = 32'h0;
    {bank3[2933], bank2[2933], bank1[2933], bank0[2933]} = 32'h0;
    {bank3[2934], bank2[2934], bank1[2934], bank0[2934]} = 32'h0;
    {bank3[2935], bank2[2935], bank1[2935], bank0[2935]} = 32'h0;
    {bank3[2936], bank2[2936], bank1[2936], bank0[2936]} = 32'h0;
    {bank3[2937], bank2[2937], bank1[2937], bank0[2937]} = 32'h0;
    {bank3[2938], bank2[2938], bank1[2938], bank0[2938]} = 32'h0;
    {bank3[2939], bank2[2939], bank1[2939], bank0[2939]} = 32'h0;
    {bank3[2940], bank2[2940], bank1[2940], bank0[2940]} = 32'h0;
    {bank3[2941], bank2[2941], bank1[2941], bank0[2941]} = 32'h0;
    {bank3[2942], bank2[2942], bank1[2942], bank0[2942]} = 32'h0;
    {bank3[2943], bank2[2943], bank1[2943], bank0[2943]} = 32'h0;
    {bank3[2944], bank2[2944], bank1[2944], bank0[2944]} = 32'h0;
    {bank3[2945], bank2[2945], bank1[2945], bank0[2945]} = 32'h0;
    {bank3[2946], bank2[2946], bank1[2946], bank0[2946]} = 32'h0;
    {bank3[2947], bank2[2947], bank1[2947], bank0[2947]} = 32'h0;
    {bank3[2948], bank2[2948], bank1[2948], bank0[2948]} = 32'h0;
    {bank3[2949], bank2[2949], bank1[2949], bank0[2949]} = 32'h0;
    {bank3[2950], bank2[2950], bank1[2950], bank0[2950]} = 32'h0;
    {bank3[2951], bank2[2951], bank1[2951], bank0[2951]} = 32'h0;
    {bank3[2952], bank2[2952], bank1[2952], bank0[2952]} = 32'h0;
    {bank3[2953], bank2[2953], bank1[2953], bank0[2953]} = 32'h0;
    {bank3[2954], bank2[2954], bank1[2954], bank0[2954]} = 32'h0;
    {bank3[2955], bank2[2955], bank1[2955], bank0[2955]} = 32'h0;
    {bank3[2956], bank2[2956], bank1[2956], bank0[2956]} = 32'h0;
    {bank3[2957], bank2[2957], bank1[2957], bank0[2957]} = 32'h0;
    {bank3[2958], bank2[2958], bank1[2958], bank0[2958]} = 32'h0;
    {bank3[2959], bank2[2959], bank1[2959], bank0[2959]} = 32'h0;
    {bank3[2960], bank2[2960], bank1[2960], bank0[2960]} = 32'h0;
    {bank3[2961], bank2[2961], bank1[2961], bank0[2961]} = 32'h0;
    {bank3[2962], bank2[2962], bank1[2962], bank0[2962]} = 32'h0;
    {bank3[2963], bank2[2963], bank1[2963], bank0[2963]} = 32'h0;
    {bank3[2964], bank2[2964], bank1[2964], bank0[2964]} = 32'h0;
    {bank3[2965], bank2[2965], bank1[2965], bank0[2965]} = 32'h0;
    {bank3[2966], bank2[2966], bank1[2966], bank0[2966]} = 32'h0;
    {bank3[2967], bank2[2967], bank1[2967], bank0[2967]} = 32'h0;
    {bank3[2968], bank2[2968], bank1[2968], bank0[2968]} = 32'h0;
    {bank3[2969], bank2[2969], bank1[2969], bank0[2969]} = 32'h0;
    {bank3[2970], bank2[2970], bank1[2970], bank0[2970]} = 32'h0;
    {bank3[2971], bank2[2971], bank1[2971], bank0[2971]} = 32'h0;
    {bank3[2972], bank2[2972], bank1[2972], bank0[2972]} = 32'h0;
    {bank3[2973], bank2[2973], bank1[2973], bank0[2973]} = 32'h0;
    {bank3[2974], bank2[2974], bank1[2974], bank0[2974]} = 32'h0;
    {bank3[2975], bank2[2975], bank1[2975], bank0[2975]} = 32'h0;
    {bank3[2976], bank2[2976], bank1[2976], bank0[2976]} = 32'h0;
    {bank3[2977], bank2[2977], bank1[2977], bank0[2977]} = 32'h0;
    {bank3[2978], bank2[2978], bank1[2978], bank0[2978]} = 32'h0;
    {bank3[2979], bank2[2979], bank1[2979], bank0[2979]} = 32'h0;
    {bank3[2980], bank2[2980], bank1[2980], bank0[2980]} = 32'h0;
    {bank3[2981], bank2[2981], bank1[2981], bank0[2981]} = 32'h0;
    {bank3[2982], bank2[2982], bank1[2982], bank0[2982]} = 32'h0;
    {bank3[2983], bank2[2983], bank1[2983], bank0[2983]} = 32'h0;
    {bank3[2984], bank2[2984], bank1[2984], bank0[2984]} = 32'h0;
    {bank3[2985], bank2[2985], bank1[2985], bank0[2985]} = 32'h0;
    {bank3[2986], bank2[2986], bank1[2986], bank0[2986]} = 32'h0;
    {bank3[2987], bank2[2987], bank1[2987], bank0[2987]} = 32'h0;
    {bank3[2988], bank2[2988], bank1[2988], bank0[2988]} = 32'h0;
    {bank3[2989], bank2[2989], bank1[2989], bank0[2989]} = 32'h0;
    {bank3[2990], bank2[2990], bank1[2990], bank0[2990]} = 32'h0;
    {bank3[2991], bank2[2991], bank1[2991], bank0[2991]} = 32'h0;
    {bank3[2992], bank2[2992], bank1[2992], bank0[2992]} = 32'h0;
    {bank3[2993], bank2[2993], bank1[2993], bank0[2993]} = 32'h0;
    {bank3[2994], bank2[2994], bank1[2994], bank0[2994]} = 32'h0;
    {bank3[2995], bank2[2995], bank1[2995], bank0[2995]} = 32'h0;
    {bank3[2996], bank2[2996], bank1[2996], bank0[2996]} = 32'h0;
    {bank3[2997], bank2[2997], bank1[2997], bank0[2997]} = 32'h0;
    {bank3[2998], bank2[2998], bank1[2998], bank0[2998]} = 32'h0;
    {bank3[2999], bank2[2999], bank1[2999], bank0[2999]} = 32'h0;
    {bank3[3000], bank2[3000], bank1[3000], bank0[3000]} = 32'h0;
    {bank3[3001], bank2[3001], bank1[3001], bank0[3001]} = 32'h0;
    {bank3[3002], bank2[3002], bank1[3002], bank0[3002]} = 32'h0;
    {bank3[3003], bank2[3003], bank1[3003], bank0[3003]} = 32'h0;
    {bank3[3004], bank2[3004], bank1[3004], bank0[3004]} = 32'h0;
    {bank3[3005], bank2[3005], bank1[3005], bank0[3005]} = 32'h0;
    {bank3[3006], bank2[3006], bank1[3006], bank0[3006]} = 32'h0;
    {bank3[3007], bank2[3007], bank1[3007], bank0[3007]} = 32'h0;
    {bank3[3008], bank2[3008], bank1[3008], bank0[3008]} = 32'h0;
    {bank3[3009], bank2[3009], bank1[3009], bank0[3009]} = 32'h0;
    {bank3[3010], bank2[3010], bank1[3010], bank0[3010]} = 32'h0;
    {bank3[3011], bank2[3011], bank1[3011], bank0[3011]} = 32'h0;
    {bank3[3012], bank2[3012], bank1[3012], bank0[3012]} = 32'h0;
    {bank3[3013], bank2[3013], bank1[3013], bank0[3013]} = 32'h0;
    {bank3[3014], bank2[3014], bank1[3014], bank0[3014]} = 32'h0;
    {bank3[3015], bank2[3015], bank1[3015], bank0[3015]} = 32'h0;
    {bank3[3016], bank2[3016], bank1[3016], bank0[3016]} = 32'h0;
    {bank3[3017], bank2[3017], bank1[3017], bank0[3017]} = 32'h0;
    {bank3[3018], bank2[3018], bank1[3018], bank0[3018]} = 32'h0;
    {bank3[3019], bank2[3019], bank1[3019], bank0[3019]} = 32'h0;
    {bank3[3020], bank2[3020], bank1[3020], bank0[3020]} = 32'h0;
    {bank3[3021], bank2[3021], bank1[3021], bank0[3021]} = 32'h0;
    {bank3[3022], bank2[3022], bank1[3022], bank0[3022]} = 32'h0;
    {bank3[3023], bank2[3023], bank1[3023], bank0[3023]} = 32'h0;
    {bank3[3024], bank2[3024], bank1[3024], bank0[3024]} = 32'h0;
    {bank3[3025], bank2[3025], bank1[3025], bank0[3025]} = 32'h0;
    {bank3[3026], bank2[3026], bank1[3026], bank0[3026]} = 32'h0;
    {bank3[3027], bank2[3027], bank1[3027], bank0[3027]} = 32'h0;
    {bank3[3028], bank2[3028], bank1[3028], bank0[3028]} = 32'h0;
    {bank3[3029], bank2[3029], bank1[3029], bank0[3029]} = 32'h0;
    {bank3[3030], bank2[3030], bank1[3030], bank0[3030]} = 32'h0;
    {bank3[3031], bank2[3031], bank1[3031], bank0[3031]} = 32'h0;
    {bank3[3032], bank2[3032], bank1[3032], bank0[3032]} = 32'h0;
    {bank3[3033], bank2[3033], bank1[3033], bank0[3033]} = 32'h0;
    {bank3[3034], bank2[3034], bank1[3034], bank0[3034]} = 32'h0;
    {bank3[3035], bank2[3035], bank1[3035], bank0[3035]} = 32'h0;
    {bank3[3036], bank2[3036], bank1[3036], bank0[3036]} = 32'h0;
    {bank3[3037], bank2[3037], bank1[3037], bank0[3037]} = 32'h0;
    {bank3[3038], bank2[3038], bank1[3038], bank0[3038]} = 32'h0;
    {bank3[3039], bank2[3039], bank1[3039], bank0[3039]} = 32'h0;
    {bank3[3040], bank2[3040], bank1[3040], bank0[3040]} = 32'h0;
    {bank3[3041], bank2[3041], bank1[3041], bank0[3041]} = 32'h0;
    {bank3[3042], bank2[3042], bank1[3042], bank0[3042]} = 32'h0;
    {bank3[3043], bank2[3043], bank1[3043], bank0[3043]} = 32'h0;
    {bank3[3044], bank2[3044], bank1[3044], bank0[3044]} = 32'h0;
    {bank3[3045], bank2[3045], bank1[3045], bank0[3045]} = 32'h0;
    {bank3[3046], bank2[3046], bank1[3046], bank0[3046]} = 32'h0;
    {bank3[3047], bank2[3047], bank1[3047], bank0[3047]} = 32'h0;
    {bank3[3048], bank2[3048], bank1[3048], bank0[3048]} = 32'h0;
    {bank3[3049], bank2[3049], bank1[3049], bank0[3049]} = 32'h0;
    {bank3[3050], bank2[3050], bank1[3050], bank0[3050]} = 32'h0;
    {bank3[3051], bank2[3051], bank1[3051], bank0[3051]} = 32'h0;
    {bank3[3052], bank2[3052], bank1[3052], bank0[3052]} = 32'h0;
    {bank3[3053], bank2[3053], bank1[3053], bank0[3053]} = 32'h0;
    {bank3[3054], bank2[3054], bank1[3054], bank0[3054]} = 32'h0;
    {bank3[3055], bank2[3055], bank1[3055], bank0[3055]} = 32'h0;
    {bank3[3056], bank2[3056], bank1[3056], bank0[3056]} = 32'h0;
    {bank3[3057], bank2[3057], bank1[3057], bank0[3057]} = 32'h0;
    {bank3[3058], bank2[3058], bank1[3058], bank0[3058]} = 32'h0;
    {bank3[3059], bank2[3059], bank1[3059], bank0[3059]} = 32'h0;
    {bank3[3060], bank2[3060], bank1[3060], bank0[3060]} = 32'h0;
    {bank3[3061], bank2[3061], bank1[3061], bank0[3061]} = 32'h0;
    {bank3[3062], bank2[3062], bank1[3062], bank0[3062]} = 32'h0;
    {bank3[3063], bank2[3063], bank1[3063], bank0[3063]} = 32'h0;
    {bank3[3064], bank2[3064], bank1[3064], bank0[3064]} = 32'h0;
    {bank3[3065], bank2[3065], bank1[3065], bank0[3065]} = 32'h0;
    {bank3[3066], bank2[3066], bank1[3066], bank0[3066]} = 32'h0;
    {bank3[3067], bank2[3067], bank1[3067], bank0[3067]} = 32'h0;
    {bank3[3068], bank2[3068], bank1[3068], bank0[3068]} = 32'h0;
    {bank3[3069], bank2[3069], bank1[3069], bank0[3069]} = 32'h0;
    {bank3[3070], bank2[3070], bank1[3070], bank0[3070]} = 32'h0;
    {bank3[3071], bank2[3071], bank1[3071], bank0[3071]} = 32'h0;
    {bank3[3072], bank2[3072], bank1[3072], bank0[3072]} = 32'h0;
    {bank3[3073], bank2[3073], bank1[3073], bank0[3073]} = 32'h0;
    {bank3[3074], bank2[3074], bank1[3074], bank0[3074]} = 32'h0;
    {bank3[3075], bank2[3075], bank1[3075], bank0[3075]} = 32'h0;
    {bank3[3076], bank2[3076], bank1[3076], bank0[3076]} = 32'h0;
    {bank3[3077], bank2[3077], bank1[3077], bank0[3077]} = 32'h0;
    {bank3[3078], bank2[3078], bank1[3078], bank0[3078]} = 32'h0;
    {bank3[3079], bank2[3079], bank1[3079], bank0[3079]} = 32'h0;
    {bank3[3080], bank2[3080], bank1[3080], bank0[3080]} = 32'h0;
    {bank3[3081], bank2[3081], bank1[3081], bank0[3081]} = 32'h0;
    {bank3[3082], bank2[3082], bank1[3082], bank0[3082]} = 32'h0;
    {bank3[3083], bank2[3083], bank1[3083], bank0[3083]} = 32'h0;
    {bank3[3084], bank2[3084], bank1[3084], bank0[3084]} = 32'h0;
    {bank3[3085], bank2[3085], bank1[3085], bank0[3085]} = 32'h0;
    {bank3[3086], bank2[3086], bank1[3086], bank0[3086]} = 32'h0;
    {bank3[3087], bank2[3087], bank1[3087], bank0[3087]} = 32'h0;
    {bank3[3088], bank2[3088], bank1[3088], bank0[3088]} = 32'h0;
    {bank3[3089], bank2[3089], bank1[3089], bank0[3089]} = 32'h0;
    {bank3[3090], bank2[3090], bank1[3090], bank0[3090]} = 32'h0;
    {bank3[3091], bank2[3091], bank1[3091], bank0[3091]} = 32'h0;
    {bank3[3092], bank2[3092], bank1[3092], bank0[3092]} = 32'h0;
    {bank3[3093], bank2[3093], bank1[3093], bank0[3093]} = 32'h0;
    {bank3[3094], bank2[3094], bank1[3094], bank0[3094]} = 32'h0;
    {bank3[3095], bank2[3095], bank1[3095], bank0[3095]} = 32'h0;
    {bank3[3096], bank2[3096], bank1[3096], bank0[3096]} = 32'h0;
    {bank3[3097], bank2[3097], bank1[3097], bank0[3097]} = 32'h0;
    {bank3[3098], bank2[3098], bank1[3098], bank0[3098]} = 32'h0;
    {bank3[3099], bank2[3099], bank1[3099], bank0[3099]} = 32'h0;
    {bank3[3100], bank2[3100], bank1[3100], bank0[3100]} = 32'h0;
    {bank3[3101], bank2[3101], bank1[3101], bank0[3101]} = 32'h0;
    {bank3[3102], bank2[3102], bank1[3102], bank0[3102]} = 32'h0;
    {bank3[3103], bank2[3103], bank1[3103], bank0[3103]} = 32'h0;
    {bank3[3104], bank2[3104], bank1[3104], bank0[3104]} = 32'h0;
    {bank3[3105], bank2[3105], bank1[3105], bank0[3105]} = 32'h0;
    {bank3[3106], bank2[3106], bank1[3106], bank0[3106]} = 32'h0;
    {bank3[3107], bank2[3107], bank1[3107], bank0[3107]} = 32'h0;
    {bank3[3108], bank2[3108], bank1[3108], bank0[3108]} = 32'h0;
    {bank3[3109], bank2[3109], bank1[3109], bank0[3109]} = 32'h0;
    {bank3[3110], bank2[3110], bank1[3110], bank0[3110]} = 32'h0;
    {bank3[3111], bank2[3111], bank1[3111], bank0[3111]} = 32'h0;
    {bank3[3112], bank2[3112], bank1[3112], bank0[3112]} = 32'h0;
    {bank3[3113], bank2[3113], bank1[3113], bank0[3113]} = 32'h0;
    {bank3[3114], bank2[3114], bank1[3114], bank0[3114]} = 32'h0;
    {bank3[3115], bank2[3115], bank1[3115], bank0[3115]} = 32'h0;
    {bank3[3116], bank2[3116], bank1[3116], bank0[3116]} = 32'h0;
    {bank3[3117], bank2[3117], bank1[3117], bank0[3117]} = 32'h0;
    {bank3[3118], bank2[3118], bank1[3118], bank0[3118]} = 32'h0;
    {bank3[3119], bank2[3119], bank1[3119], bank0[3119]} = 32'h0;
    {bank3[3120], bank2[3120], bank1[3120], bank0[3120]} = 32'h0;
    {bank3[3121], bank2[3121], bank1[3121], bank0[3121]} = 32'h0;
    {bank3[3122], bank2[3122], bank1[3122], bank0[3122]} = 32'h0;
    {bank3[3123], bank2[3123], bank1[3123], bank0[3123]} = 32'h0;
    {bank3[3124], bank2[3124], bank1[3124], bank0[3124]} = 32'h0;
    {bank3[3125], bank2[3125], bank1[3125], bank0[3125]} = 32'h0;
    {bank3[3126], bank2[3126], bank1[3126], bank0[3126]} = 32'h0;
    {bank3[3127], bank2[3127], bank1[3127], bank0[3127]} = 32'h0;
    {bank3[3128], bank2[3128], bank1[3128], bank0[3128]} = 32'h0;
    {bank3[3129], bank2[3129], bank1[3129], bank0[3129]} = 32'h0;
    {bank3[3130], bank2[3130], bank1[3130], bank0[3130]} = 32'h0;
    {bank3[3131], bank2[3131], bank1[3131], bank0[3131]} = 32'h0;
    {bank3[3132], bank2[3132], bank1[3132], bank0[3132]} = 32'h0;
    {bank3[3133], bank2[3133], bank1[3133], bank0[3133]} = 32'h0;
    {bank3[3134], bank2[3134], bank1[3134], bank0[3134]} = 32'h0;
    {bank3[3135], bank2[3135], bank1[3135], bank0[3135]} = 32'h0;
    {bank3[3136], bank2[3136], bank1[3136], bank0[3136]} = 32'h0;
    {bank3[3137], bank2[3137], bank1[3137], bank0[3137]} = 32'h0;
    {bank3[3138], bank2[3138], bank1[3138], bank0[3138]} = 32'h0;
    {bank3[3139], bank2[3139], bank1[3139], bank0[3139]} = 32'h0;
    {bank3[3140], bank2[3140], bank1[3140], bank0[3140]} = 32'h0;
    {bank3[3141], bank2[3141], bank1[3141], bank0[3141]} = 32'h0;
    {bank3[3142], bank2[3142], bank1[3142], bank0[3142]} = 32'h0;
    {bank3[3143], bank2[3143], bank1[3143], bank0[3143]} = 32'h0;
    {bank3[3144], bank2[3144], bank1[3144], bank0[3144]} = 32'h0;
    {bank3[3145], bank2[3145], bank1[3145], bank0[3145]} = 32'h0;
    {bank3[3146], bank2[3146], bank1[3146], bank0[3146]} = 32'h0;
    {bank3[3147], bank2[3147], bank1[3147], bank0[3147]} = 32'h0;
    {bank3[3148], bank2[3148], bank1[3148], bank0[3148]} = 32'h0;
    {bank3[3149], bank2[3149], bank1[3149], bank0[3149]} = 32'h0;
    {bank3[3150], bank2[3150], bank1[3150], bank0[3150]} = 32'h0;
    {bank3[3151], bank2[3151], bank1[3151], bank0[3151]} = 32'h0;
    {bank3[3152], bank2[3152], bank1[3152], bank0[3152]} = 32'h0;
    {bank3[3153], bank2[3153], bank1[3153], bank0[3153]} = 32'h0;
    {bank3[3154], bank2[3154], bank1[3154], bank0[3154]} = 32'h0;
    {bank3[3155], bank2[3155], bank1[3155], bank0[3155]} = 32'h0;
    {bank3[3156], bank2[3156], bank1[3156], bank0[3156]} = 32'h0;
    {bank3[3157], bank2[3157], bank1[3157], bank0[3157]} = 32'h0;
    {bank3[3158], bank2[3158], bank1[3158], bank0[3158]} = 32'h0;
    {bank3[3159], bank2[3159], bank1[3159], bank0[3159]} = 32'h0;
    {bank3[3160], bank2[3160], bank1[3160], bank0[3160]} = 32'h0;
    {bank3[3161], bank2[3161], bank1[3161], bank0[3161]} = 32'h0;
    {bank3[3162], bank2[3162], bank1[3162], bank0[3162]} = 32'h0;
    {bank3[3163], bank2[3163], bank1[3163], bank0[3163]} = 32'h0;
    {bank3[3164], bank2[3164], bank1[3164], bank0[3164]} = 32'h0;
    {bank3[3165], bank2[3165], bank1[3165], bank0[3165]} = 32'h0;
    {bank3[3166], bank2[3166], bank1[3166], bank0[3166]} = 32'h0;
    {bank3[3167], bank2[3167], bank1[3167], bank0[3167]} = 32'h0;
    {bank3[3168], bank2[3168], bank1[3168], bank0[3168]} = 32'h0;
    {bank3[3169], bank2[3169], bank1[3169], bank0[3169]} = 32'h0;
    {bank3[3170], bank2[3170], bank1[3170], bank0[3170]} = 32'h0;
    {bank3[3171], bank2[3171], bank1[3171], bank0[3171]} = 32'h0;
    {bank3[3172], bank2[3172], bank1[3172], bank0[3172]} = 32'h0;
    {bank3[3173], bank2[3173], bank1[3173], bank0[3173]} = 32'h0;
    {bank3[3174], bank2[3174], bank1[3174], bank0[3174]} = 32'h0;
    {bank3[3175], bank2[3175], bank1[3175], bank0[3175]} = 32'h0;
    {bank3[3176], bank2[3176], bank1[3176], bank0[3176]} = 32'h0;
    {bank3[3177], bank2[3177], bank1[3177], bank0[3177]} = 32'h0;
    {bank3[3178], bank2[3178], bank1[3178], bank0[3178]} = 32'h0;
    {bank3[3179], bank2[3179], bank1[3179], bank0[3179]} = 32'h0;
    {bank3[3180], bank2[3180], bank1[3180], bank0[3180]} = 32'h0;
    {bank3[3181], bank2[3181], bank1[3181], bank0[3181]} = 32'h0;
    {bank3[3182], bank2[3182], bank1[3182], bank0[3182]} = 32'h0;
    {bank3[3183], bank2[3183], bank1[3183], bank0[3183]} = 32'h0;
    {bank3[3184], bank2[3184], bank1[3184], bank0[3184]} = 32'h0;
    {bank3[3185], bank2[3185], bank1[3185], bank0[3185]} = 32'h0;
    {bank3[3186], bank2[3186], bank1[3186], bank0[3186]} = 32'h0;
    {bank3[3187], bank2[3187], bank1[3187], bank0[3187]} = 32'h0;
    {bank3[3188], bank2[3188], bank1[3188], bank0[3188]} = 32'h0;
    {bank3[3189], bank2[3189], bank1[3189], bank0[3189]} = 32'h0;
    {bank3[3190], bank2[3190], bank1[3190], bank0[3190]} = 32'h0;
    {bank3[3191], bank2[3191], bank1[3191], bank0[3191]} = 32'h0;
    {bank3[3192], bank2[3192], bank1[3192], bank0[3192]} = 32'h0;
    {bank3[3193], bank2[3193], bank1[3193], bank0[3193]} = 32'h0;
    {bank3[3194], bank2[3194], bank1[3194], bank0[3194]} = 32'h0;
    {bank3[3195], bank2[3195], bank1[3195], bank0[3195]} = 32'h0;
    {bank3[3196], bank2[3196], bank1[3196], bank0[3196]} = 32'h0;
    {bank3[3197], bank2[3197], bank1[3197], bank0[3197]} = 32'h0;
    {bank3[3198], bank2[3198], bank1[3198], bank0[3198]} = 32'h0;
    {bank3[3199], bank2[3199], bank1[3199], bank0[3199]} = 32'h0;
    {bank3[3200], bank2[3200], bank1[3200], bank0[3200]} = 32'h0;
    {bank3[3201], bank2[3201], bank1[3201], bank0[3201]} = 32'h0;
    {bank3[3202], bank2[3202], bank1[3202], bank0[3202]} = 32'h0;
    {bank3[3203], bank2[3203], bank1[3203], bank0[3203]} = 32'h0;
    {bank3[3204], bank2[3204], bank1[3204], bank0[3204]} = 32'h0;
    {bank3[3205], bank2[3205], bank1[3205], bank0[3205]} = 32'h0;
    {bank3[3206], bank2[3206], bank1[3206], bank0[3206]} = 32'h0;
    {bank3[3207], bank2[3207], bank1[3207], bank0[3207]} = 32'h0;
    {bank3[3208], bank2[3208], bank1[3208], bank0[3208]} = 32'h0;
    {bank3[3209], bank2[3209], bank1[3209], bank0[3209]} = 32'h0;
    {bank3[3210], bank2[3210], bank1[3210], bank0[3210]} = 32'h0;
    {bank3[3211], bank2[3211], bank1[3211], bank0[3211]} = 32'h0;
    {bank3[3212], bank2[3212], bank1[3212], bank0[3212]} = 32'h0;
    {bank3[3213], bank2[3213], bank1[3213], bank0[3213]} = 32'h0;
    {bank3[3214], bank2[3214], bank1[3214], bank0[3214]} = 32'h0;
    {bank3[3215], bank2[3215], bank1[3215], bank0[3215]} = 32'h0;
    {bank3[3216], bank2[3216], bank1[3216], bank0[3216]} = 32'h0;
    {bank3[3217], bank2[3217], bank1[3217], bank0[3217]} = 32'h0;
    {bank3[3218], bank2[3218], bank1[3218], bank0[3218]} = 32'h0;
    {bank3[3219], bank2[3219], bank1[3219], bank0[3219]} = 32'h0;
    {bank3[3220], bank2[3220], bank1[3220], bank0[3220]} = 32'h0;
    {bank3[3221], bank2[3221], bank1[3221], bank0[3221]} = 32'h0;
    {bank3[3222], bank2[3222], bank1[3222], bank0[3222]} = 32'h0;
    {bank3[3223], bank2[3223], bank1[3223], bank0[3223]} = 32'h0;
    {bank3[3224], bank2[3224], bank1[3224], bank0[3224]} = 32'h0;
    {bank3[3225], bank2[3225], bank1[3225], bank0[3225]} = 32'h0;
    {bank3[3226], bank2[3226], bank1[3226], bank0[3226]} = 32'h0;
    {bank3[3227], bank2[3227], bank1[3227], bank0[3227]} = 32'h0;
    {bank3[3228], bank2[3228], bank1[3228], bank0[3228]} = 32'h0;
    {bank3[3229], bank2[3229], bank1[3229], bank0[3229]} = 32'h0;
    {bank3[3230], bank2[3230], bank1[3230], bank0[3230]} = 32'h0;
    {bank3[3231], bank2[3231], bank1[3231], bank0[3231]} = 32'h0;
    {bank3[3232], bank2[3232], bank1[3232], bank0[3232]} = 32'h0;
    {bank3[3233], bank2[3233], bank1[3233], bank0[3233]} = 32'h0;
    {bank3[3234], bank2[3234], bank1[3234], bank0[3234]} = 32'h0;
    {bank3[3235], bank2[3235], bank1[3235], bank0[3235]} = 32'h0;
    {bank3[3236], bank2[3236], bank1[3236], bank0[3236]} = 32'h0;
    {bank3[3237], bank2[3237], bank1[3237], bank0[3237]} = 32'h0;
    {bank3[3238], bank2[3238], bank1[3238], bank0[3238]} = 32'h0;
    {bank3[3239], bank2[3239], bank1[3239], bank0[3239]} = 32'h0;
    {bank3[3240], bank2[3240], bank1[3240], bank0[3240]} = 32'h0;
    {bank3[3241], bank2[3241], bank1[3241], bank0[3241]} = 32'h0;
    {bank3[3242], bank2[3242], bank1[3242], bank0[3242]} = 32'h0;
    {bank3[3243], bank2[3243], bank1[3243], bank0[3243]} = 32'h0;
    {bank3[3244], bank2[3244], bank1[3244], bank0[3244]} = 32'h0;
    {bank3[3245], bank2[3245], bank1[3245], bank0[3245]} = 32'h0;
    {bank3[3246], bank2[3246], bank1[3246], bank0[3246]} = 32'h0;
    {bank3[3247], bank2[3247], bank1[3247], bank0[3247]} = 32'h0;
    {bank3[3248], bank2[3248], bank1[3248], bank0[3248]} = 32'h0;
    {bank3[3249], bank2[3249], bank1[3249], bank0[3249]} = 32'h0;
    {bank3[3250], bank2[3250], bank1[3250], bank0[3250]} = 32'h0;
    {bank3[3251], bank2[3251], bank1[3251], bank0[3251]} = 32'h0;
    {bank3[3252], bank2[3252], bank1[3252], bank0[3252]} = 32'h0;
    {bank3[3253], bank2[3253], bank1[3253], bank0[3253]} = 32'h0;
    {bank3[3254], bank2[3254], bank1[3254], bank0[3254]} = 32'h0;
    {bank3[3255], bank2[3255], bank1[3255], bank0[3255]} = 32'h0;
    {bank3[3256], bank2[3256], bank1[3256], bank0[3256]} = 32'h0;
    {bank3[3257], bank2[3257], bank1[3257], bank0[3257]} = 32'h0;
    {bank3[3258], bank2[3258], bank1[3258], bank0[3258]} = 32'h0;
    {bank3[3259], bank2[3259], bank1[3259], bank0[3259]} = 32'h0;
    {bank3[3260], bank2[3260], bank1[3260], bank0[3260]} = 32'h0;
    {bank3[3261], bank2[3261], bank1[3261], bank0[3261]} = 32'h0;
    {bank3[3262], bank2[3262], bank1[3262], bank0[3262]} = 32'h0;
    {bank3[3263], bank2[3263], bank1[3263], bank0[3263]} = 32'h0;
    {bank3[3264], bank2[3264], bank1[3264], bank0[3264]} = 32'h0;
    {bank3[3265], bank2[3265], bank1[3265], bank0[3265]} = 32'h0;
    {bank3[3266], bank2[3266], bank1[3266], bank0[3266]} = 32'h0;
    {bank3[3267], bank2[3267], bank1[3267], bank0[3267]} = 32'h0;
    {bank3[3268], bank2[3268], bank1[3268], bank0[3268]} = 32'h0;
    {bank3[3269], bank2[3269], bank1[3269], bank0[3269]} = 32'h0;
    {bank3[3270], bank2[3270], bank1[3270], bank0[3270]} = 32'h0;
    {bank3[3271], bank2[3271], bank1[3271], bank0[3271]} = 32'h0;
    {bank3[3272], bank2[3272], bank1[3272], bank0[3272]} = 32'h0;
    {bank3[3273], bank2[3273], bank1[3273], bank0[3273]} = 32'h0;
    {bank3[3274], bank2[3274], bank1[3274], bank0[3274]} = 32'h0;
    {bank3[3275], bank2[3275], bank1[3275], bank0[3275]} = 32'h0;
    {bank3[3276], bank2[3276], bank1[3276], bank0[3276]} = 32'h0;
    {bank3[3277], bank2[3277], bank1[3277], bank0[3277]} = 32'h0;
    {bank3[3278], bank2[3278], bank1[3278], bank0[3278]} = 32'h0;
    {bank3[3279], bank2[3279], bank1[3279], bank0[3279]} = 32'h0;
    {bank3[3280], bank2[3280], bank1[3280], bank0[3280]} = 32'h0;
    {bank3[3281], bank2[3281], bank1[3281], bank0[3281]} = 32'h0;
    {bank3[3282], bank2[3282], bank1[3282], bank0[3282]} = 32'h0;
    {bank3[3283], bank2[3283], bank1[3283], bank0[3283]} = 32'h0;
    {bank3[3284], bank2[3284], bank1[3284], bank0[3284]} = 32'h0;
    {bank3[3285], bank2[3285], bank1[3285], bank0[3285]} = 32'h0;
    {bank3[3286], bank2[3286], bank1[3286], bank0[3286]} = 32'h0;
    {bank3[3287], bank2[3287], bank1[3287], bank0[3287]} = 32'h0;
    {bank3[3288], bank2[3288], bank1[3288], bank0[3288]} = 32'h0;
    {bank3[3289], bank2[3289], bank1[3289], bank0[3289]} = 32'h0;
    {bank3[3290], bank2[3290], bank1[3290], bank0[3290]} = 32'h0;
    {bank3[3291], bank2[3291], bank1[3291], bank0[3291]} = 32'h0;
    {bank3[3292], bank2[3292], bank1[3292], bank0[3292]} = 32'h0;
    {bank3[3293], bank2[3293], bank1[3293], bank0[3293]} = 32'h0;
    {bank3[3294], bank2[3294], bank1[3294], bank0[3294]} = 32'h0;
    {bank3[3295], bank2[3295], bank1[3295], bank0[3295]} = 32'h0;
    {bank3[3296], bank2[3296], bank1[3296], bank0[3296]} = 32'h0;
    {bank3[3297], bank2[3297], bank1[3297], bank0[3297]} = 32'h0;
    {bank3[3298], bank2[3298], bank1[3298], bank0[3298]} = 32'h0;
    {bank3[3299], bank2[3299], bank1[3299], bank0[3299]} = 32'h0;
    {bank3[3300], bank2[3300], bank1[3300], bank0[3300]} = 32'h0;
    {bank3[3301], bank2[3301], bank1[3301], bank0[3301]} = 32'h0;
    {bank3[3302], bank2[3302], bank1[3302], bank0[3302]} = 32'h0;
    {bank3[3303], bank2[3303], bank1[3303], bank0[3303]} = 32'h0;
    {bank3[3304], bank2[3304], bank1[3304], bank0[3304]} = 32'h0;
    {bank3[3305], bank2[3305], bank1[3305], bank0[3305]} = 32'h0;
    {bank3[3306], bank2[3306], bank1[3306], bank0[3306]} = 32'h0;
    {bank3[3307], bank2[3307], bank1[3307], bank0[3307]} = 32'h0;
    {bank3[3308], bank2[3308], bank1[3308], bank0[3308]} = 32'h0;
    {bank3[3309], bank2[3309], bank1[3309], bank0[3309]} = 32'h0;
    {bank3[3310], bank2[3310], bank1[3310], bank0[3310]} = 32'h0;
    {bank3[3311], bank2[3311], bank1[3311], bank0[3311]} = 32'h0;
    {bank3[3312], bank2[3312], bank1[3312], bank0[3312]} = 32'h0;
    {bank3[3313], bank2[3313], bank1[3313], bank0[3313]} = 32'h0;
    {bank3[3314], bank2[3314], bank1[3314], bank0[3314]} = 32'h0;
    {bank3[3315], bank2[3315], bank1[3315], bank0[3315]} = 32'h0;
    {bank3[3316], bank2[3316], bank1[3316], bank0[3316]} = 32'h0;
    {bank3[3317], bank2[3317], bank1[3317], bank0[3317]} = 32'h0;
    {bank3[3318], bank2[3318], bank1[3318], bank0[3318]} = 32'h0;
    {bank3[3319], bank2[3319], bank1[3319], bank0[3319]} = 32'h0;
    {bank3[3320], bank2[3320], bank1[3320], bank0[3320]} = 32'h0;
    {bank3[3321], bank2[3321], bank1[3321], bank0[3321]} = 32'h0;
    {bank3[3322], bank2[3322], bank1[3322], bank0[3322]} = 32'h0;
    {bank3[3323], bank2[3323], bank1[3323], bank0[3323]} = 32'h0;
    {bank3[3324], bank2[3324], bank1[3324], bank0[3324]} = 32'h0;
    {bank3[3325], bank2[3325], bank1[3325], bank0[3325]} = 32'h0;
    {bank3[3326], bank2[3326], bank1[3326], bank0[3326]} = 32'h0;
    {bank3[3327], bank2[3327], bank1[3327], bank0[3327]} = 32'h0;
    {bank3[3328], bank2[3328], bank1[3328], bank0[3328]} = 32'h0;
    {bank3[3329], bank2[3329], bank1[3329], bank0[3329]} = 32'h0;
    {bank3[3330], bank2[3330], bank1[3330], bank0[3330]} = 32'h0;
    {bank3[3331], bank2[3331], bank1[3331], bank0[3331]} = 32'h0;
    {bank3[3332], bank2[3332], bank1[3332], bank0[3332]} = 32'h0;
    {bank3[3333], bank2[3333], bank1[3333], bank0[3333]} = 32'h0;
    {bank3[3334], bank2[3334], bank1[3334], bank0[3334]} = 32'h0;
    {bank3[3335], bank2[3335], bank1[3335], bank0[3335]} = 32'h0;
    {bank3[3336], bank2[3336], bank1[3336], bank0[3336]} = 32'h0;
    {bank3[3337], bank2[3337], bank1[3337], bank0[3337]} = 32'h0;
    {bank3[3338], bank2[3338], bank1[3338], bank0[3338]} = 32'h0;
    {bank3[3339], bank2[3339], bank1[3339], bank0[3339]} = 32'h0;
    {bank3[3340], bank2[3340], bank1[3340], bank0[3340]} = 32'h0;
    {bank3[3341], bank2[3341], bank1[3341], bank0[3341]} = 32'h0;
    {bank3[3342], bank2[3342], bank1[3342], bank0[3342]} = 32'h0;
    {bank3[3343], bank2[3343], bank1[3343], bank0[3343]} = 32'h0;
    {bank3[3344], bank2[3344], bank1[3344], bank0[3344]} = 32'h0;
    {bank3[3345], bank2[3345], bank1[3345], bank0[3345]} = 32'h0;
    {bank3[3346], bank2[3346], bank1[3346], bank0[3346]} = 32'h0;
    {bank3[3347], bank2[3347], bank1[3347], bank0[3347]} = 32'h0;
    {bank3[3348], bank2[3348], bank1[3348], bank0[3348]} = 32'h0;
    {bank3[3349], bank2[3349], bank1[3349], bank0[3349]} = 32'h0;
    {bank3[3350], bank2[3350], bank1[3350], bank0[3350]} = 32'h0;
    {bank3[3351], bank2[3351], bank1[3351], bank0[3351]} = 32'h0;
    {bank3[3352], bank2[3352], bank1[3352], bank0[3352]} = 32'h0;
    {bank3[3353], bank2[3353], bank1[3353], bank0[3353]} = 32'h0;
    {bank3[3354], bank2[3354], bank1[3354], bank0[3354]} = 32'h0;
    {bank3[3355], bank2[3355], bank1[3355], bank0[3355]} = 32'h0;
    {bank3[3356], bank2[3356], bank1[3356], bank0[3356]} = 32'h0;
    {bank3[3357], bank2[3357], bank1[3357], bank0[3357]} = 32'h0;
    {bank3[3358], bank2[3358], bank1[3358], bank0[3358]} = 32'h0;
    {bank3[3359], bank2[3359], bank1[3359], bank0[3359]} = 32'h0;
    {bank3[3360], bank2[3360], bank1[3360], bank0[3360]} = 32'h0;
    {bank3[3361], bank2[3361], bank1[3361], bank0[3361]} = 32'h0;
    {bank3[3362], bank2[3362], bank1[3362], bank0[3362]} = 32'h0;
    {bank3[3363], bank2[3363], bank1[3363], bank0[3363]} = 32'h0;
    {bank3[3364], bank2[3364], bank1[3364], bank0[3364]} = 32'h0;
    {bank3[3365], bank2[3365], bank1[3365], bank0[3365]} = 32'h0;
    {bank3[3366], bank2[3366], bank1[3366], bank0[3366]} = 32'h0;
    {bank3[3367], bank2[3367], bank1[3367], bank0[3367]} = 32'h0;
    {bank3[3368], bank2[3368], bank1[3368], bank0[3368]} = 32'h0;
    {bank3[3369], bank2[3369], bank1[3369], bank0[3369]} = 32'h0;
    {bank3[3370], bank2[3370], bank1[3370], bank0[3370]} = 32'h0;
    {bank3[3371], bank2[3371], bank1[3371], bank0[3371]} = 32'h0;
    {bank3[3372], bank2[3372], bank1[3372], bank0[3372]} = 32'h0;
    {bank3[3373], bank2[3373], bank1[3373], bank0[3373]} = 32'h0;
    {bank3[3374], bank2[3374], bank1[3374], bank0[3374]} = 32'h0;
    {bank3[3375], bank2[3375], bank1[3375], bank0[3375]} = 32'h0;
    {bank3[3376], bank2[3376], bank1[3376], bank0[3376]} = 32'h0;
    {bank3[3377], bank2[3377], bank1[3377], bank0[3377]} = 32'h0;
    {bank3[3378], bank2[3378], bank1[3378], bank0[3378]} = 32'h0;
    {bank3[3379], bank2[3379], bank1[3379], bank0[3379]} = 32'h0;
    {bank3[3380], bank2[3380], bank1[3380], bank0[3380]} = 32'h0;
    {bank3[3381], bank2[3381], bank1[3381], bank0[3381]} = 32'h0;
    {bank3[3382], bank2[3382], bank1[3382], bank0[3382]} = 32'h0;
    {bank3[3383], bank2[3383], bank1[3383], bank0[3383]} = 32'h0;
    {bank3[3384], bank2[3384], bank1[3384], bank0[3384]} = 32'h0;
    {bank3[3385], bank2[3385], bank1[3385], bank0[3385]} = 32'h0;
    {bank3[3386], bank2[3386], bank1[3386], bank0[3386]} = 32'h0;
    {bank3[3387], bank2[3387], bank1[3387], bank0[3387]} = 32'h0;
    {bank3[3388], bank2[3388], bank1[3388], bank0[3388]} = 32'h0;
    {bank3[3389], bank2[3389], bank1[3389], bank0[3389]} = 32'h0;
    {bank3[3390], bank2[3390], bank1[3390], bank0[3390]} = 32'h0;
    {bank3[3391], bank2[3391], bank1[3391], bank0[3391]} = 32'h0;
    {bank3[3392], bank2[3392], bank1[3392], bank0[3392]} = 32'h0;
    {bank3[3393], bank2[3393], bank1[3393], bank0[3393]} = 32'h0;
    {bank3[3394], bank2[3394], bank1[3394], bank0[3394]} = 32'h0;
    {bank3[3395], bank2[3395], bank1[3395], bank0[3395]} = 32'h0;
    {bank3[3396], bank2[3396], bank1[3396], bank0[3396]} = 32'h0;
    {bank3[3397], bank2[3397], bank1[3397], bank0[3397]} = 32'h0;
    {bank3[3398], bank2[3398], bank1[3398], bank0[3398]} = 32'h0;
    {bank3[3399], bank2[3399], bank1[3399], bank0[3399]} = 32'h0;
    {bank3[3400], bank2[3400], bank1[3400], bank0[3400]} = 32'h0;
    {bank3[3401], bank2[3401], bank1[3401], bank0[3401]} = 32'h0;
    {bank3[3402], bank2[3402], bank1[3402], bank0[3402]} = 32'h0;
    {bank3[3403], bank2[3403], bank1[3403], bank0[3403]} = 32'h0;
    {bank3[3404], bank2[3404], bank1[3404], bank0[3404]} = 32'h0;
    {bank3[3405], bank2[3405], bank1[3405], bank0[3405]} = 32'h0;
    {bank3[3406], bank2[3406], bank1[3406], bank0[3406]} = 32'h0;
    {bank3[3407], bank2[3407], bank1[3407], bank0[3407]} = 32'h0;
    {bank3[3408], bank2[3408], bank1[3408], bank0[3408]} = 32'h0;
    {bank3[3409], bank2[3409], bank1[3409], bank0[3409]} = 32'h0;
    {bank3[3410], bank2[3410], bank1[3410], bank0[3410]} = 32'h0;
    {bank3[3411], bank2[3411], bank1[3411], bank0[3411]} = 32'h0;
    {bank3[3412], bank2[3412], bank1[3412], bank0[3412]} = 32'h0;
    {bank3[3413], bank2[3413], bank1[3413], bank0[3413]} = 32'h0;
    {bank3[3414], bank2[3414], bank1[3414], bank0[3414]} = 32'h0;
    {bank3[3415], bank2[3415], bank1[3415], bank0[3415]} = 32'h0;
    {bank3[3416], bank2[3416], bank1[3416], bank0[3416]} = 32'h0;
    {bank3[3417], bank2[3417], bank1[3417], bank0[3417]} = 32'h0;
    {bank3[3418], bank2[3418], bank1[3418], bank0[3418]} = 32'h0;
    {bank3[3419], bank2[3419], bank1[3419], bank0[3419]} = 32'h0;
    {bank3[3420], bank2[3420], bank1[3420], bank0[3420]} = 32'h0;
    {bank3[3421], bank2[3421], bank1[3421], bank0[3421]} = 32'h0;
    {bank3[3422], bank2[3422], bank1[3422], bank0[3422]} = 32'h0;
    {bank3[3423], bank2[3423], bank1[3423], bank0[3423]} = 32'h0;
    {bank3[3424], bank2[3424], bank1[3424], bank0[3424]} = 32'h0;
    {bank3[3425], bank2[3425], bank1[3425], bank0[3425]} = 32'h0;
    {bank3[3426], bank2[3426], bank1[3426], bank0[3426]} = 32'h0;
    {bank3[3427], bank2[3427], bank1[3427], bank0[3427]} = 32'h0;
    {bank3[3428], bank2[3428], bank1[3428], bank0[3428]} = 32'h0;
    {bank3[3429], bank2[3429], bank1[3429], bank0[3429]} = 32'h0;
    {bank3[3430], bank2[3430], bank1[3430], bank0[3430]} = 32'h0;
    {bank3[3431], bank2[3431], bank1[3431], bank0[3431]} = 32'h0;
    {bank3[3432], bank2[3432], bank1[3432], bank0[3432]} = 32'h0;
    {bank3[3433], bank2[3433], bank1[3433], bank0[3433]} = 32'h0;
    {bank3[3434], bank2[3434], bank1[3434], bank0[3434]} = 32'h0;
    {bank3[3435], bank2[3435], bank1[3435], bank0[3435]} = 32'h0;
    {bank3[3436], bank2[3436], bank1[3436], bank0[3436]} = 32'h0;
    {bank3[3437], bank2[3437], bank1[3437], bank0[3437]} = 32'h0;
    {bank3[3438], bank2[3438], bank1[3438], bank0[3438]} = 32'h0;
    {bank3[3439], bank2[3439], bank1[3439], bank0[3439]} = 32'h0;
    {bank3[3440], bank2[3440], bank1[3440], bank0[3440]} = 32'h0;
    {bank3[3441], bank2[3441], bank1[3441], bank0[3441]} = 32'h0;
    {bank3[3442], bank2[3442], bank1[3442], bank0[3442]} = 32'h0;
    {bank3[3443], bank2[3443], bank1[3443], bank0[3443]} = 32'h0;
    {bank3[3444], bank2[3444], bank1[3444], bank0[3444]} = 32'h0;
    {bank3[3445], bank2[3445], bank1[3445], bank0[3445]} = 32'h0;
    {bank3[3446], bank2[3446], bank1[3446], bank0[3446]} = 32'h0;
    {bank3[3447], bank2[3447], bank1[3447], bank0[3447]} = 32'h0;
    {bank3[3448], bank2[3448], bank1[3448], bank0[3448]} = 32'h0;
    {bank3[3449], bank2[3449], bank1[3449], bank0[3449]} = 32'h0;
    {bank3[3450], bank2[3450], bank1[3450], bank0[3450]} = 32'h0;
    {bank3[3451], bank2[3451], bank1[3451], bank0[3451]} = 32'h0;
    {bank3[3452], bank2[3452], bank1[3452], bank0[3452]} = 32'h0;
    {bank3[3453], bank2[3453], bank1[3453], bank0[3453]} = 32'h0;
    {bank3[3454], bank2[3454], bank1[3454], bank0[3454]} = 32'h0;
    {bank3[3455], bank2[3455], bank1[3455], bank0[3455]} = 32'h0;
    {bank3[3456], bank2[3456], bank1[3456], bank0[3456]} = 32'h0;
    {bank3[3457], bank2[3457], bank1[3457], bank0[3457]} = 32'h0;
    {bank3[3458], bank2[3458], bank1[3458], bank0[3458]} = 32'h0;
    {bank3[3459], bank2[3459], bank1[3459], bank0[3459]} = 32'h0;
    {bank3[3460], bank2[3460], bank1[3460], bank0[3460]} = 32'h0;
    {bank3[3461], bank2[3461], bank1[3461], bank0[3461]} = 32'h0;
    {bank3[3462], bank2[3462], bank1[3462], bank0[3462]} = 32'h0;
    {bank3[3463], bank2[3463], bank1[3463], bank0[3463]} = 32'h0;
    {bank3[3464], bank2[3464], bank1[3464], bank0[3464]} = 32'h0;
    {bank3[3465], bank2[3465], bank1[3465], bank0[3465]} = 32'h0;
    {bank3[3466], bank2[3466], bank1[3466], bank0[3466]} = 32'h0;
    {bank3[3467], bank2[3467], bank1[3467], bank0[3467]} = 32'h0;
    {bank3[3468], bank2[3468], bank1[3468], bank0[3468]} = 32'h0;
    {bank3[3469], bank2[3469], bank1[3469], bank0[3469]} = 32'h0;
    {bank3[3470], bank2[3470], bank1[3470], bank0[3470]} = 32'h0;
    {bank3[3471], bank2[3471], bank1[3471], bank0[3471]} = 32'h0;
    {bank3[3472], bank2[3472], bank1[3472], bank0[3472]} = 32'h0;
    {bank3[3473], bank2[3473], bank1[3473], bank0[3473]} = 32'h0;
    {bank3[3474], bank2[3474], bank1[3474], bank0[3474]} = 32'h0;
    {bank3[3475], bank2[3475], bank1[3475], bank0[3475]} = 32'h0;
    {bank3[3476], bank2[3476], bank1[3476], bank0[3476]} = 32'h0;
    {bank3[3477], bank2[3477], bank1[3477], bank0[3477]} = 32'h0;
    {bank3[3478], bank2[3478], bank1[3478], bank0[3478]} = 32'h0;
    {bank3[3479], bank2[3479], bank1[3479], bank0[3479]} = 32'h0;
    {bank3[3480], bank2[3480], bank1[3480], bank0[3480]} = 32'h0;
    {bank3[3481], bank2[3481], bank1[3481], bank0[3481]} = 32'h0;
    {bank3[3482], bank2[3482], bank1[3482], bank0[3482]} = 32'h0;
    {bank3[3483], bank2[3483], bank1[3483], bank0[3483]} = 32'h0;
    {bank3[3484], bank2[3484], bank1[3484], bank0[3484]} = 32'h0;
    {bank3[3485], bank2[3485], bank1[3485], bank0[3485]} = 32'h0;
    {bank3[3486], bank2[3486], bank1[3486], bank0[3486]} = 32'h0;
    {bank3[3487], bank2[3487], bank1[3487], bank0[3487]} = 32'h0;
    {bank3[3488], bank2[3488], bank1[3488], bank0[3488]} = 32'h0;
    {bank3[3489], bank2[3489], bank1[3489], bank0[3489]} = 32'h0;
    {bank3[3490], bank2[3490], bank1[3490], bank0[3490]} = 32'h0;
    {bank3[3491], bank2[3491], bank1[3491], bank0[3491]} = 32'h0;
    {bank3[3492], bank2[3492], bank1[3492], bank0[3492]} = 32'h0;
    {bank3[3493], bank2[3493], bank1[3493], bank0[3493]} = 32'h0;
    {bank3[3494], bank2[3494], bank1[3494], bank0[3494]} = 32'h0;
    {bank3[3495], bank2[3495], bank1[3495], bank0[3495]} = 32'h0;
    {bank3[3496], bank2[3496], bank1[3496], bank0[3496]} = 32'h0;
    {bank3[3497], bank2[3497], bank1[3497], bank0[3497]} = 32'h0;
    {bank3[3498], bank2[3498], bank1[3498], bank0[3498]} = 32'h0;
    {bank3[3499], bank2[3499], bank1[3499], bank0[3499]} = 32'h0;
    {bank3[3500], bank2[3500], bank1[3500], bank0[3500]} = 32'h0;
    {bank3[3501], bank2[3501], bank1[3501], bank0[3501]} = 32'h0;
    {bank3[3502], bank2[3502], bank1[3502], bank0[3502]} = 32'h0;
    {bank3[3503], bank2[3503], bank1[3503], bank0[3503]} = 32'h0;
    {bank3[3504], bank2[3504], bank1[3504], bank0[3504]} = 32'h0;
    {bank3[3505], bank2[3505], bank1[3505], bank0[3505]} = 32'h0;
    {bank3[3506], bank2[3506], bank1[3506], bank0[3506]} = 32'h0;
    {bank3[3507], bank2[3507], bank1[3507], bank0[3507]} = 32'h0;
    {bank3[3508], bank2[3508], bank1[3508], bank0[3508]} = 32'h0;
    {bank3[3509], bank2[3509], bank1[3509], bank0[3509]} = 32'h0;
    {bank3[3510], bank2[3510], bank1[3510], bank0[3510]} = 32'h0;
    {bank3[3511], bank2[3511], bank1[3511], bank0[3511]} = 32'h0;
    {bank3[3512], bank2[3512], bank1[3512], bank0[3512]} = 32'h0;
    {bank3[3513], bank2[3513], bank1[3513], bank0[3513]} = 32'h0;
    {bank3[3514], bank2[3514], bank1[3514], bank0[3514]} = 32'h0;
    {bank3[3515], bank2[3515], bank1[3515], bank0[3515]} = 32'h0;
    {bank3[3516], bank2[3516], bank1[3516], bank0[3516]} = 32'h0;
    {bank3[3517], bank2[3517], bank1[3517], bank0[3517]} = 32'h0;
    {bank3[3518], bank2[3518], bank1[3518], bank0[3518]} = 32'h0;
    {bank3[3519], bank2[3519], bank1[3519], bank0[3519]} = 32'h0;
    {bank3[3520], bank2[3520], bank1[3520], bank0[3520]} = 32'h0;
    {bank3[3521], bank2[3521], bank1[3521], bank0[3521]} = 32'h0;
    {bank3[3522], bank2[3522], bank1[3522], bank0[3522]} = 32'h0;
    {bank3[3523], bank2[3523], bank1[3523], bank0[3523]} = 32'h0;
    {bank3[3524], bank2[3524], bank1[3524], bank0[3524]} = 32'h0;
    {bank3[3525], bank2[3525], bank1[3525], bank0[3525]} = 32'h0;
    {bank3[3526], bank2[3526], bank1[3526], bank0[3526]} = 32'h0;
    {bank3[3527], bank2[3527], bank1[3527], bank0[3527]} = 32'h0;
    {bank3[3528], bank2[3528], bank1[3528], bank0[3528]} = 32'h0;
    {bank3[3529], bank2[3529], bank1[3529], bank0[3529]} = 32'h0;
    {bank3[3530], bank2[3530], bank1[3530], bank0[3530]} = 32'h0;
    {bank3[3531], bank2[3531], bank1[3531], bank0[3531]} = 32'h0;
    {bank3[3532], bank2[3532], bank1[3532], bank0[3532]} = 32'h0;
    {bank3[3533], bank2[3533], bank1[3533], bank0[3533]} = 32'h0;
    {bank3[3534], bank2[3534], bank1[3534], bank0[3534]} = 32'h0;
    {bank3[3535], bank2[3535], bank1[3535], bank0[3535]} = 32'h0;
    {bank3[3536], bank2[3536], bank1[3536], bank0[3536]} = 32'h0;
    {bank3[3537], bank2[3537], bank1[3537], bank0[3537]} = 32'h0;
    {bank3[3538], bank2[3538], bank1[3538], bank0[3538]} = 32'h0;
    {bank3[3539], bank2[3539], bank1[3539], bank0[3539]} = 32'h0;
    {bank3[3540], bank2[3540], bank1[3540], bank0[3540]} = 32'h0;
    {bank3[3541], bank2[3541], bank1[3541], bank0[3541]} = 32'h0;
    {bank3[3542], bank2[3542], bank1[3542], bank0[3542]} = 32'h0;
    {bank3[3543], bank2[3543], bank1[3543], bank0[3543]} = 32'h0;
    {bank3[3544], bank2[3544], bank1[3544], bank0[3544]} = 32'h0;
    {bank3[3545], bank2[3545], bank1[3545], bank0[3545]} = 32'h0;
    {bank3[3546], bank2[3546], bank1[3546], bank0[3546]} = 32'h0;
    {bank3[3547], bank2[3547], bank1[3547], bank0[3547]} = 32'h0;
    {bank3[3548], bank2[3548], bank1[3548], bank0[3548]} = 32'h0;
    {bank3[3549], bank2[3549], bank1[3549], bank0[3549]} = 32'h0;
    {bank3[3550], bank2[3550], bank1[3550], bank0[3550]} = 32'h0;
    {bank3[3551], bank2[3551], bank1[3551], bank0[3551]} = 32'h0;
    {bank3[3552], bank2[3552], bank1[3552], bank0[3552]} = 32'h0;
    {bank3[3553], bank2[3553], bank1[3553], bank0[3553]} = 32'h0;
    {bank3[3554], bank2[3554], bank1[3554], bank0[3554]} = 32'h0;
    {bank3[3555], bank2[3555], bank1[3555], bank0[3555]} = 32'h0;
    {bank3[3556], bank2[3556], bank1[3556], bank0[3556]} = 32'h0;
    {bank3[3557], bank2[3557], bank1[3557], bank0[3557]} = 32'h0;
    {bank3[3558], bank2[3558], bank1[3558], bank0[3558]} = 32'h0;
    {bank3[3559], bank2[3559], bank1[3559], bank0[3559]} = 32'h0;
    {bank3[3560], bank2[3560], bank1[3560], bank0[3560]} = 32'h0;
    {bank3[3561], bank2[3561], bank1[3561], bank0[3561]} = 32'h0;
    {bank3[3562], bank2[3562], bank1[3562], bank0[3562]} = 32'h0;
    {bank3[3563], bank2[3563], bank1[3563], bank0[3563]} = 32'h0;
    {bank3[3564], bank2[3564], bank1[3564], bank0[3564]} = 32'h0;
    {bank3[3565], bank2[3565], bank1[3565], bank0[3565]} = 32'h0;
    {bank3[3566], bank2[3566], bank1[3566], bank0[3566]} = 32'h0;
    {bank3[3567], bank2[3567], bank1[3567], bank0[3567]} = 32'h0;
    {bank3[3568], bank2[3568], bank1[3568], bank0[3568]} = 32'h0;
    {bank3[3569], bank2[3569], bank1[3569], bank0[3569]} = 32'h0;
    {bank3[3570], bank2[3570], bank1[3570], bank0[3570]} = 32'h0;
    {bank3[3571], bank2[3571], bank1[3571], bank0[3571]} = 32'h0;
    {bank3[3572], bank2[3572], bank1[3572], bank0[3572]} = 32'h0;
    {bank3[3573], bank2[3573], bank1[3573], bank0[3573]} = 32'h0;
    {bank3[3574], bank2[3574], bank1[3574], bank0[3574]} = 32'h0;
    {bank3[3575], bank2[3575], bank1[3575], bank0[3575]} = 32'h0;
    {bank3[3576], bank2[3576], bank1[3576], bank0[3576]} = 32'h0;
    {bank3[3577], bank2[3577], bank1[3577], bank0[3577]} = 32'h0;
    {bank3[3578], bank2[3578], bank1[3578], bank0[3578]} = 32'h0;
    {bank3[3579], bank2[3579], bank1[3579], bank0[3579]} = 32'h0;
    {bank3[3580], bank2[3580], bank1[3580], bank0[3580]} = 32'h0;
    {bank3[3581], bank2[3581], bank1[3581], bank0[3581]} = 32'h0;
    {bank3[3582], bank2[3582], bank1[3582], bank0[3582]} = 32'h0;
    {bank3[3583], bank2[3583], bank1[3583], bank0[3583]} = 32'h0;
    {bank3[3584], bank2[3584], bank1[3584], bank0[3584]} = 32'h0;
    {bank3[3585], bank2[3585], bank1[3585], bank0[3585]} = 32'h0;
    {bank3[3586], bank2[3586], bank1[3586], bank0[3586]} = 32'h0;
    {bank3[3587], bank2[3587], bank1[3587], bank0[3587]} = 32'h0;
    {bank3[3588], bank2[3588], bank1[3588], bank0[3588]} = 32'h0;
    {bank3[3589], bank2[3589], bank1[3589], bank0[3589]} = 32'h0;
    {bank3[3590], bank2[3590], bank1[3590], bank0[3590]} = 32'h0;
    {bank3[3591], bank2[3591], bank1[3591], bank0[3591]} = 32'h0;
    {bank3[3592], bank2[3592], bank1[3592], bank0[3592]} = 32'h0;
    {bank3[3593], bank2[3593], bank1[3593], bank0[3593]} = 32'h0;
    {bank3[3594], bank2[3594], bank1[3594], bank0[3594]} = 32'h0;
    {bank3[3595], bank2[3595], bank1[3595], bank0[3595]} = 32'h0;
    {bank3[3596], bank2[3596], bank1[3596], bank0[3596]} = 32'h0;
    {bank3[3597], bank2[3597], bank1[3597], bank0[3597]} = 32'h0;
    {bank3[3598], bank2[3598], bank1[3598], bank0[3598]} = 32'h0;
    {bank3[3599], bank2[3599], bank1[3599], bank0[3599]} = 32'h0;
    {bank3[3600], bank2[3600], bank1[3600], bank0[3600]} = 32'h0;
    {bank3[3601], bank2[3601], bank1[3601], bank0[3601]} = 32'h0;
    {bank3[3602], bank2[3602], bank1[3602], bank0[3602]} = 32'h0;
    {bank3[3603], bank2[3603], bank1[3603], bank0[3603]} = 32'h0;
    {bank3[3604], bank2[3604], bank1[3604], bank0[3604]} = 32'h0;
    {bank3[3605], bank2[3605], bank1[3605], bank0[3605]} = 32'h0;
    {bank3[3606], bank2[3606], bank1[3606], bank0[3606]} = 32'h0;
    {bank3[3607], bank2[3607], bank1[3607], bank0[3607]} = 32'h0;
    {bank3[3608], bank2[3608], bank1[3608], bank0[3608]} = 32'h0;
    {bank3[3609], bank2[3609], bank1[3609], bank0[3609]} = 32'h0;
    {bank3[3610], bank2[3610], bank1[3610], bank0[3610]} = 32'h0;
    {bank3[3611], bank2[3611], bank1[3611], bank0[3611]} = 32'h0;
    {bank3[3612], bank2[3612], bank1[3612], bank0[3612]} = 32'h0;
    {bank3[3613], bank2[3613], bank1[3613], bank0[3613]} = 32'h0;
    {bank3[3614], bank2[3614], bank1[3614], bank0[3614]} = 32'h0;
    {bank3[3615], bank2[3615], bank1[3615], bank0[3615]} = 32'h0;
    {bank3[3616], bank2[3616], bank1[3616], bank0[3616]} = 32'h0;
    {bank3[3617], bank2[3617], bank1[3617], bank0[3617]} = 32'h0;
    {bank3[3618], bank2[3618], bank1[3618], bank0[3618]} = 32'h0;
    {bank3[3619], bank2[3619], bank1[3619], bank0[3619]} = 32'h0;
    {bank3[3620], bank2[3620], bank1[3620], bank0[3620]} = 32'h0;
    {bank3[3621], bank2[3621], bank1[3621], bank0[3621]} = 32'h0;
    {bank3[3622], bank2[3622], bank1[3622], bank0[3622]} = 32'h0;
    {bank3[3623], bank2[3623], bank1[3623], bank0[3623]} = 32'h0;
    {bank3[3624], bank2[3624], bank1[3624], bank0[3624]} = 32'h0;
    {bank3[3625], bank2[3625], bank1[3625], bank0[3625]} = 32'h0;
    {bank3[3626], bank2[3626], bank1[3626], bank0[3626]} = 32'h0;
    {bank3[3627], bank2[3627], bank1[3627], bank0[3627]} = 32'h0;
    {bank3[3628], bank2[3628], bank1[3628], bank0[3628]} = 32'h0;
    {bank3[3629], bank2[3629], bank1[3629], bank0[3629]} = 32'h0;
    {bank3[3630], bank2[3630], bank1[3630], bank0[3630]} = 32'h0;
    {bank3[3631], bank2[3631], bank1[3631], bank0[3631]} = 32'h0;
    {bank3[3632], bank2[3632], bank1[3632], bank0[3632]} = 32'h0;
    {bank3[3633], bank2[3633], bank1[3633], bank0[3633]} = 32'h0;
    {bank3[3634], bank2[3634], bank1[3634], bank0[3634]} = 32'h0;
    {bank3[3635], bank2[3635], bank1[3635], bank0[3635]} = 32'h0;
    {bank3[3636], bank2[3636], bank1[3636], bank0[3636]} = 32'h0;
    {bank3[3637], bank2[3637], bank1[3637], bank0[3637]} = 32'h0;
    {bank3[3638], bank2[3638], bank1[3638], bank0[3638]} = 32'h0;
    {bank3[3639], bank2[3639], bank1[3639], bank0[3639]} = 32'h0;
    {bank3[3640], bank2[3640], bank1[3640], bank0[3640]} = 32'h0;
    {bank3[3641], bank2[3641], bank1[3641], bank0[3641]} = 32'h0;
    {bank3[3642], bank2[3642], bank1[3642], bank0[3642]} = 32'h0;
    {bank3[3643], bank2[3643], bank1[3643], bank0[3643]} = 32'h0;
    {bank3[3644], bank2[3644], bank1[3644], bank0[3644]} = 32'h0;
    {bank3[3645], bank2[3645], bank1[3645], bank0[3645]} = 32'h0;
    {bank3[3646], bank2[3646], bank1[3646], bank0[3646]} = 32'h0;
    {bank3[3647], bank2[3647], bank1[3647], bank0[3647]} = 32'h0;
    {bank3[3648], bank2[3648], bank1[3648], bank0[3648]} = 32'h0;
    {bank3[3649], bank2[3649], bank1[3649], bank0[3649]} = 32'h0;
    {bank3[3650], bank2[3650], bank1[3650], bank0[3650]} = 32'h0;
    {bank3[3651], bank2[3651], bank1[3651], bank0[3651]} = 32'h0;
    {bank3[3652], bank2[3652], bank1[3652], bank0[3652]} = 32'h0;
    {bank3[3653], bank2[3653], bank1[3653], bank0[3653]} = 32'h0;
    {bank3[3654], bank2[3654], bank1[3654], bank0[3654]} = 32'h0;
    {bank3[3655], bank2[3655], bank1[3655], bank0[3655]} = 32'h0;
    {bank3[3656], bank2[3656], bank1[3656], bank0[3656]} = 32'h0;
    {bank3[3657], bank2[3657], bank1[3657], bank0[3657]} = 32'h0;
    {bank3[3658], bank2[3658], bank1[3658], bank0[3658]} = 32'h0;
    {bank3[3659], bank2[3659], bank1[3659], bank0[3659]} = 32'h0;
    {bank3[3660], bank2[3660], bank1[3660], bank0[3660]} = 32'h0;
    {bank3[3661], bank2[3661], bank1[3661], bank0[3661]} = 32'h0;
    {bank3[3662], bank2[3662], bank1[3662], bank0[3662]} = 32'h0;
    {bank3[3663], bank2[3663], bank1[3663], bank0[3663]} = 32'h0;
    {bank3[3664], bank2[3664], bank1[3664], bank0[3664]} = 32'h0;
    {bank3[3665], bank2[3665], bank1[3665], bank0[3665]} = 32'h0;
    {bank3[3666], bank2[3666], bank1[3666], bank0[3666]} = 32'h0;
    {bank3[3667], bank2[3667], bank1[3667], bank0[3667]} = 32'h0;
    {bank3[3668], bank2[3668], bank1[3668], bank0[3668]} = 32'h0;
    {bank3[3669], bank2[3669], bank1[3669], bank0[3669]} = 32'h0;
    {bank3[3670], bank2[3670], bank1[3670], bank0[3670]} = 32'h0;
    {bank3[3671], bank2[3671], bank1[3671], bank0[3671]} = 32'h0;
    {bank3[3672], bank2[3672], bank1[3672], bank0[3672]} = 32'h0;
    {bank3[3673], bank2[3673], bank1[3673], bank0[3673]} = 32'h0;
    {bank3[3674], bank2[3674], bank1[3674], bank0[3674]} = 32'h0;
    {bank3[3675], bank2[3675], bank1[3675], bank0[3675]} = 32'h0;
    {bank3[3676], bank2[3676], bank1[3676], bank0[3676]} = 32'h0;
    {bank3[3677], bank2[3677], bank1[3677], bank0[3677]} = 32'h0;
    {bank3[3678], bank2[3678], bank1[3678], bank0[3678]} = 32'h0;
    {bank3[3679], bank2[3679], bank1[3679], bank0[3679]} = 32'h0;
    {bank3[3680], bank2[3680], bank1[3680], bank0[3680]} = 32'h0;
    {bank3[3681], bank2[3681], bank1[3681], bank0[3681]} = 32'h0;
    {bank3[3682], bank2[3682], bank1[3682], bank0[3682]} = 32'h0;
    {bank3[3683], bank2[3683], bank1[3683], bank0[3683]} = 32'h0;
    {bank3[3684], bank2[3684], bank1[3684], bank0[3684]} = 32'h0;
    {bank3[3685], bank2[3685], bank1[3685], bank0[3685]} = 32'h0;
    {bank3[3686], bank2[3686], bank1[3686], bank0[3686]} = 32'h0;
    {bank3[3687], bank2[3687], bank1[3687], bank0[3687]} = 32'h0;
    {bank3[3688], bank2[3688], bank1[3688], bank0[3688]} = 32'h0;
    {bank3[3689], bank2[3689], bank1[3689], bank0[3689]} = 32'h0;
    {bank3[3690], bank2[3690], bank1[3690], bank0[3690]} = 32'h0;
    {bank3[3691], bank2[3691], bank1[3691], bank0[3691]} = 32'h0;
    {bank3[3692], bank2[3692], bank1[3692], bank0[3692]} = 32'h0;
    {bank3[3693], bank2[3693], bank1[3693], bank0[3693]} = 32'h0;
    {bank3[3694], bank2[3694], bank1[3694], bank0[3694]} = 32'h0;
    {bank3[3695], bank2[3695], bank1[3695], bank0[3695]} = 32'h0;
    {bank3[3696], bank2[3696], bank1[3696], bank0[3696]} = 32'h0;
    {bank3[3697], bank2[3697], bank1[3697], bank0[3697]} = 32'h0;
    {bank3[3698], bank2[3698], bank1[3698], bank0[3698]} = 32'h0;
    {bank3[3699], bank2[3699], bank1[3699], bank0[3699]} = 32'h0;
    {bank3[3700], bank2[3700], bank1[3700], bank0[3700]} = 32'h0;
    {bank3[3701], bank2[3701], bank1[3701], bank0[3701]} = 32'h0;
    {bank3[3702], bank2[3702], bank1[3702], bank0[3702]} = 32'h0;
    {bank3[3703], bank2[3703], bank1[3703], bank0[3703]} = 32'h0;
    {bank3[3704], bank2[3704], bank1[3704], bank0[3704]} = 32'h0;
    {bank3[3705], bank2[3705], bank1[3705], bank0[3705]} = 32'h0;
    {bank3[3706], bank2[3706], bank1[3706], bank0[3706]} = 32'h0;
    {bank3[3707], bank2[3707], bank1[3707], bank0[3707]} = 32'h0;
    {bank3[3708], bank2[3708], bank1[3708], bank0[3708]} = 32'h0;
    {bank3[3709], bank2[3709], bank1[3709], bank0[3709]} = 32'h0;
    {bank3[3710], bank2[3710], bank1[3710], bank0[3710]} = 32'h0;
    {bank3[3711], bank2[3711], bank1[3711], bank0[3711]} = 32'h0;
    {bank3[3712], bank2[3712], bank1[3712], bank0[3712]} = 32'h0;
    {bank3[3713], bank2[3713], bank1[3713], bank0[3713]} = 32'h0;
    {bank3[3714], bank2[3714], bank1[3714], bank0[3714]} = 32'h0;
    {bank3[3715], bank2[3715], bank1[3715], bank0[3715]} = 32'h0;
    {bank3[3716], bank2[3716], bank1[3716], bank0[3716]} = 32'h0;
    {bank3[3717], bank2[3717], bank1[3717], bank0[3717]} = 32'h0;
    {bank3[3718], bank2[3718], bank1[3718], bank0[3718]} = 32'h0;
    {bank3[3719], bank2[3719], bank1[3719], bank0[3719]} = 32'h0;
    {bank3[3720], bank2[3720], bank1[3720], bank0[3720]} = 32'h0;
    {bank3[3721], bank2[3721], bank1[3721], bank0[3721]} = 32'h0;
    {bank3[3722], bank2[3722], bank1[3722], bank0[3722]} = 32'h0;
    {bank3[3723], bank2[3723], bank1[3723], bank0[3723]} = 32'h0;
    {bank3[3724], bank2[3724], bank1[3724], bank0[3724]} = 32'h0;
    {bank3[3725], bank2[3725], bank1[3725], bank0[3725]} = 32'h0;
    {bank3[3726], bank2[3726], bank1[3726], bank0[3726]} = 32'h0;
    {bank3[3727], bank2[3727], bank1[3727], bank0[3727]} = 32'h0;
    {bank3[3728], bank2[3728], bank1[3728], bank0[3728]} = 32'h0;
    {bank3[3729], bank2[3729], bank1[3729], bank0[3729]} = 32'h0;
    {bank3[3730], bank2[3730], bank1[3730], bank0[3730]} = 32'h0;
    {bank3[3731], bank2[3731], bank1[3731], bank0[3731]} = 32'h0;
    {bank3[3732], bank2[3732], bank1[3732], bank0[3732]} = 32'h0;
    {bank3[3733], bank2[3733], bank1[3733], bank0[3733]} = 32'h0;
    {bank3[3734], bank2[3734], bank1[3734], bank0[3734]} = 32'h0;
    {bank3[3735], bank2[3735], bank1[3735], bank0[3735]} = 32'h0;
    {bank3[3736], bank2[3736], bank1[3736], bank0[3736]} = 32'h0;
    {bank3[3737], bank2[3737], bank1[3737], bank0[3737]} = 32'h0;
    {bank3[3738], bank2[3738], bank1[3738], bank0[3738]} = 32'h0;
    {bank3[3739], bank2[3739], bank1[3739], bank0[3739]} = 32'h0;
    {bank3[3740], bank2[3740], bank1[3740], bank0[3740]} = 32'h0;
    {bank3[3741], bank2[3741], bank1[3741], bank0[3741]} = 32'h0;
    {bank3[3742], bank2[3742], bank1[3742], bank0[3742]} = 32'h0;
    {bank3[3743], bank2[3743], bank1[3743], bank0[3743]} = 32'h0;
    {bank3[3744], bank2[3744], bank1[3744], bank0[3744]} = 32'h0;
    {bank3[3745], bank2[3745], bank1[3745], bank0[3745]} = 32'h0;
    {bank3[3746], bank2[3746], bank1[3746], bank0[3746]} = 32'h0;
    {bank3[3747], bank2[3747], bank1[3747], bank0[3747]} = 32'h0;
    {bank3[3748], bank2[3748], bank1[3748], bank0[3748]} = 32'h0;
    {bank3[3749], bank2[3749], bank1[3749], bank0[3749]} = 32'h0;
    {bank3[3750], bank2[3750], bank1[3750], bank0[3750]} = 32'h0;
    {bank3[3751], bank2[3751], bank1[3751], bank0[3751]} = 32'h0;
    {bank3[3752], bank2[3752], bank1[3752], bank0[3752]} = 32'h0;
    {bank3[3753], bank2[3753], bank1[3753], bank0[3753]} = 32'h0;
    {bank3[3754], bank2[3754], bank1[3754], bank0[3754]} = 32'h0;
    {bank3[3755], bank2[3755], bank1[3755], bank0[3755]} = 32'h0;
    {bank3[3756], bank2[3756], bank1[3756], bank0[3756]} = 32'h0;
    {bank3[3757], bank2[3757], bank1[3757], bank0[3757]} = 32'h0;
    {bank3[3758], bank2[3758], bank1[3758], bank0[3758]} = 32'h0;
    {bank3[3759], bank2[3759], bank1[3759], bank0[3759]} = 32'h0;
    {bank3[3760], bank2[3760], bank1[3760], bank0[3760]} = 32'h0;
    {bank3[3761], bank2[3761], bank1[3761], bank0[3761]} = 32'h0;
    {bank3[3762], bank2[3762], bank1[3762], bank0[3762]} = 32'h0;
    {bank3[3763], bank2[3763], bank1[3763], bank0[3763]} = 32'h0;
    {bank3[3764], bank2[3764], bank1[3764], bank0[3764]} = 32'h0;
    {bank3[3765], bank2[3765], bank1[3765], bank0[3765]} = 32'h0;
    {bank3[3766], bank2[3766], bank1[3766], bank0[3766]} = 32'h0;
    {bank3[3767], bank2[3767], bank1[3767], bank0[3767]} = 32'h0;
    {bank3[3768], bank2[3768], bank1[3768], bank0[3768]} = 32'h0;
    {bank3[3769], bank2[3769], bank1[3769], bank0[3769]} = 32'h0;
    {bank3[3770], bank2[3770], bank1[3770], bank0[3770]} = 32'h0;
    {bank3[3771], bank2[3771], bank1[3771], bank0[3771]} = 32'h0;
    {bank3[3772], bank2[3772], bank1[3772], bank0[3772]} = 32'h0;
    {bank3[3773], bank2[3773], bank1[3773], bank0[3773]} = 32'h0;
    {bank3[3774], bank2[3774], bank1[3774], bank0[3774]} = 32'h0;
    {bank3[3775], bank2[3775], bank1[3775], bank0[3775]} = 32'h0;
    {bank3[3776], bank2[3776], bank1[3776], bank0[3776]} = 32'h0;
    {bank3[3777], bank2[3777], bank1[3777], bank0[3777]} = 32'h0;
    {bank3[3778], bank2[3778], bank1[3778], bank0[3778]} = 32'h0;
    {bank3[3779], bank2[3779], bank1[3779], bank0[3779]} = 32'h0;
    {bank3[3780], bank2[3780], bank1[3780], bank0[3780]} = 32'h0;
    {bank3[3781], bank2[3781], bank1[3781], bank0[3781]} = 32'h0;
    {bank3[3782], bank2[3782], bank1[3782], bank0[3782]} = 32'h0;
    {bank3[3783], bank2[3783], bank1[3783], bank0[3783]} = 32'h0;
    {bank3[3784], bank2[3784], bank1[3784], bank0[3784]} = 32'h0;
    {bank3[3785], bank2[3785], bank1[3785], bank0[3785]} = 32'h0;
    {bank3[3786], bank2[3786], bank1[3786], bank0[3786]} = 32'h0;
    {bank3[3787], bank2[3787], bank1[3787], bank0[3787]} = 32'h0;
    {bank3[3788], bank2[3788], bank1[3788], bank0[3788]} = 32'h0;
    {bank3[3789], bank2[3789], bank1[3789], bank0[3789]} = 32'h0;
    {bank3[3790], bank2[3790], bank1[3790], bank0[3790]} = 32'h0;
    {bank3[3791], bank2[3791], bank1[3791], bank0[3791]} = 32'h0;
    {bank3[3792], bank2[3792], bank1[3792], bank0[3792]} = 32'h0;
    {bank3[3793], bank2[3793], bank1[3793], bank0[3793]} = 32'h0;
    {bank3[3794], bank2[3794], bank1[3794], bank0[3794]} = 32'h0;
    {bank3[3795], bank2[3795], bank1[3795], bank0[3795]} = 32'h0;
    {bank3[3796], bank2[3796], bank1[3796], bank0[3796]} = 32'h0;
    {bank3[3797], bank2[3797], bank1[3797], bank0[3797]} = 32'h0;
    {bank3[3798], bank2[3798], bank1[3798], bank0[3798]} = 32'h0;
    {bank3[3799], bank2[3799], bank1[3799], bank0[3799]} = 32'h0;
    {bank3[3800], bank2[3800], bank1[3800], bank0[3800]} = 32'h0;
    {bank3[3801], bank2[3801], bank1[3801], bank0[3801]} = 32'h0;
    {bank3[3802], bank2[3802], bank1[3802], bank0[3802]} = 32'h0;
    {bank3[3803], bank2[3803], bank1[3803], bank0[3803]} = 32'h0;
    {bank3[3804], bank2[3804], bank1[3804], bank0[3804]} = 32'h0;
    {bank3[3805], bank2[3805], bank1[3805], bank0[3805]} = 32'h0;
    {bank3[3806], bank2[3806], bank1[3806], bank0[3806]} = 32'h0;
    {bank3[3807], bank2[3807], bank1[3807], bank0[3807]} = 32'h0;
    {bank3[3808], bank2[3808], bank1[3808], bank0[3808]} = 32'h0;
    {bank3[3809], bank2[3809], bank1[3809], bank0[3809]} = 32'h0;
    {bank3[3810], bank2[3810], bank1[3810], bank0[3810]} = 32'h0;
    {bank3[3811], bank2[3811], bank1[3811], bank0[3811]} = 32'h0;
    {bank3[3812], bank2[3812], bank1[3812], bank0[3812]} = 32'h0;
    {bank3[3813], bank2[3813], bank1[3813], bank0[3813]} = 32'h0;
    {bank3[3814], bank2[3814], bank1[3814], bank0[3814]} = 32'h0;
    {bank3[3815], bank2[3815], bank1[3815], bank0[3815]} = 32'h0;
    {bank3[3816], bank2[3816], bank1[3816], bank0[3816]} = 32'h0;
    {bank3[3817], bank2[3817], bank1[3817], bank0[3817]} = 32'h0;
    {bank3[3818], bank2[3818], bank1[3818], bank0[3818]} = 32'h0;
    {bank3[3819], bank2[3819], bank1[3819], bank0[3819]} = 32'h0;
    {bank3[3820], bank2[3820], bank1[3820], bank0[3820]} = 32'h0;
    {bank3[3821], bank2[3821], bank1[3821], bank0[3821]} = 32'h0;
    {bank3[3822], bank2[3822], bank1[3822], bank0[3822]} = 32'h0;
    {bank3[3823], bank2[3823], bank1[3823], bank0[3823]} = 32'h0;
    {bank3[3824], bank2[3824], bank1[3824], bank0[3824]} = 32'h0;
    {bank3[3825], bank2[3825], bank1[3825], bank0[3825]} = 32'h0;
    {bank3[3826], bank2[3826], bank1[3826], bank0[3826]} = 32'h0;
    {bank3[3827], bank2[3827], bank1[3827], bank0[3827]} = 32'h0;
    {bank3[3828], bank2[3828], bank1[3828], bank0[3828]} = 32'h0;
    {bank3[3829], bank2[3829], bank1[3829], bank0[3829]} = 32'h0;
    {bank3[3830], bank2[3830], bank1[3830], bank0[3830]} = 32'h0;
    {bank3[3831], bank2[3831], bank1[3831], bank0[3831]} = 32'h0;
    {bank3[3832], bank2[3832], bank1[3832], bank0[3832]} = 32'h0;
    {bank3[3833], bank2[3833], bank1[3833], bank0[3833]} = 32'h0;
    {bank3[3834], bank2[3834], bank1[3834], bank0[3834]} = 32'h0;
    {bank3[3835], bank2[3835], bank1[3835], bank0[3835]} = 32'h0;
    {bank3[3836], bank2[3836], bank1[3836], bank0[3836]} = 32'h0;
    {bank3[3837], bank2[3837], bank1[3837], bank0[3837]} = 32'h0;
    {bank3[3838], bank2[3838], bank1[3838], bank0[3838]} = 32'h0;
    {bank3[3839], bank2[3839], bank1[3839], bank0[3839]} = 32'h0;
    {bank3[3840], bank2[3840], bank1[3840], bank0[3840]} = 32'h0;
    {bank3[3841], bank2[3841], bank1[3841], bank0[3841]} = 32'h0;
    {bank3[3842], bank2[3842], bank1[3842], bank0[3842]} = 32'h0;
    {bank3[3843], bank2[3843], bank1[3843], bank0[3843]} = 32'h0;
    {bank3[3844], bank2[3844], bank1[3844], bank0[3844]} = 32'h0;
    {bank3[3845], bank2[3845], bank1[3845], bank0[3845]} = 32'h0;
    {bank3[3846], bank2[3846], bank1[3846], bank0[3846]} = 32'h0;
    {bank3[3847], bank2[3847], bank1[3847], bank0[3847]} = 32'h0;
    {bank3[3848], bank2[3848], bank1[3848], bank0[3848]} = 32'h0;
    {bank3[3849], bank2[3849], bank1[3849], bank0[3849]} = 32'h0;
    {bank3[3850], bank2[3850], bank1[3850], bank0[3850]} = 32'h0;
    {bank3[3851], bank2[3851], bank1[3851], bank0[3851]} = 32'h0;
    {bank3[3852], bank2[3852], bank1[3852], bank0[3852]} = 32'h0;
    {bank3[3853], bank2[3853], bank1[3853], bank0[3853]} = 32'h0;
    {bank3[3854], bank2[3854], bank1[3854], bank0[3854]} = 32'h0;
    {bank3[3855], bank2[3855], bank1[3855], bank0[3855]} = 32'h0;
    {bank3[3856], bank2[3856], bank1[3856], bank0[3856]} = 32'h0;
    {bank3[3857], bank2[3857], bank1[3857], bank0[3857]} = 32'h0;
    {bank3[3858], bank2[3858], bank1[3858], bank0[3858]} = 32'h0;
    {bank3[3859], bank2[3859], bank1[3859], bank0[3859]} = 32'h0;
    {bank3[3860], bank2[3860], bank1[3860], bank0[3860]} = 32'h0;
    {bank3[3861], bank2[3861], bank1[3861], bank0[3861]} = 32'h0;
    {bank3[3862], bank2[3862], bank1[3862], bank0[3862]} = 32'h0;
    {bank3[3863], bank2[3863], bank1[3863], bank0[3863]} = 32'h0;
    {bank3[3864], bank2[3864], bank1[3864], bank0[3864]} = 32'h0;
    {bank3[3865], bank2[3865], bank1[3865], bank0[3865]} = 32'h0;
    {bank3[3866], bank2[3866], bank1[3866], bank0[3866]} = 32'h0;
    {bank3[3867], bank2[3867], bank1[3867], bank0[3867]} = 32'h0;
    {bank3[3868], bank2[3868], bank1[3868], bank0[3868]} = 32'h0;
    {bank3[3869], bank2[3869], bank1[3869], bank0[3869]} = 32'h0;
    {bank3[3870], bank2[3870], bank1[3870], bank0[3870]} = 32'h0;
    {bank3[3871], bank2[3871], bank1[3871], bank0[3871]} = 32'h0;
    {bank3[3872], bank2[3872], bank1[3872], bank0[3872]} = 32'h0;
    {bank3[3873], bank2[3873], bank1[3873], bank0[3873]} = 32'h0;
    {bank3[3874], bank2[3874], bank1[3874], bank0[3874]} = 32'h0;
    {bank3[3875], bank2[3875], bank1[3875], bank0[3875]} = 32'h0;
    {bank3[3876], bank2[3876], bank1[3876], bank0[3876]} = 32'h0;
    {bank3[3877], bank2[3877], bank1[3877], bank0[3877]} = 32'h0;
    {bank3[3878], bank2[3878], bank1[3878], bank0[3878]} = 32'h0;
    {bank3[3879], bank2[3879], bank1[3879], bank0[3879]} = 32'h0;
    {bank3[3880], bank2[3880], bank1[3880], bank0[3880]} = 32'h0;
    {bank3[3881], bank2[3881], bank1[3881], bank0[3881]} = 32'h0;
    {bank3[3882], bank2[3882], bank1[3882], bank0[3882]} = 32'h0;
    {bank3[3883], bank2[3883], bank1[3883], bank0[3883]} = 32'h0;
    {bank3[3884], bank2[3884], bank1[3884], bank0[3884]} = 32'h0;
    {bank3[3885], bank2[3885], bank1[3885], bank0[3885]} = 32'h0;
    {bank3[3886], bank2[3886], bank1[3886], bank0[3886]} = 32'h0;
    {bank3[3887], bank2[3887], bank1[3887], bank0[3887]} = 32'h0;
    {bank3[3888], bank2[3888], bank1[3888], bank0[3888]} = 32'h0;
    {bank3[3889], bank2[3889], bank1[3889], bank0[3889]} = 32'h0;
    {bank3[3890], bank2[3890], bank1[3890], bank0[3890]} = 32'h0;
    {bank3[3891], bank2[3891], bank1[3891], bank0[3891]} = 32'h0;
    {bank3[3892], bank2[3892], bank1[3892], bank0[3892]} = 32'h0;
    {bank3[3893], bank2[3893], bank1[3893], bank0[3893]} = 32'h0;
    {bank3[3894], bank2[3894], bank1[3894], bank0[3894]} = 32'h0;
    {bank3[3895], bank2[3895], bank1[3895], bank0[3895]} = 32'h0;
    {bank3[3896], bank2[3896], bank1[3896], bank0[3896]} = 32'h0;
    {bank3[3897], bank2[3897], bank1[3897], bank0[3897]} = 32'h0;
    {bank3[3898], bank2[3898], bank1[3898], bank0[3898]} = 32'h0;
    {bank3[3899], bank2[3899], bank1[3899], bank0[3899]} = 32'h0;
    {bank3[3900], bank2[3900], bank1[3900], bank0[3900]} = 32'h0;
    {bank3[3901], bank2[3901], bank1[3901], bank0[3901]} = 32'h0;
    {bank3[3902], bank2[3902], bank1[3902], bank0[3902]} = 32'h0;
    {bank3[3903], bank2[3903], bank1[3903], bank0[3903]} = 32'h0;
    {bank3[3904], bank2[3904], bank1[3904], bank0[3904]} = 32'h0;
    {bank3[3905], bank2[3905], bank1[3905], bank0[3905]} = 32'h0;
    {bank3[3906], bank2[3906], bank1[3906], bank0[3906]} = 32'h0;
    {bank3[3907], bank2[3907], bank1[3907], bank0[3907]} = 32'h0;
    {bank3[3908], bank2[3908], bank1[3908], bank0[3908]} = 32'h0;
    {bank3[3909], bank2[3909], bank1[3909], bank0[3909]} = 32'h0;
    {bank3[3910], bank2[3910], bank1[3910], bank0[3910]} = 32'h0;
    {bank3[3911], bank2[3911], bank1[3911], bank0[3911]} = 32'h0;
    {bank3[3912], bank2[3912], bank1[3912], bank0[3912]} = 32'h0;
    {bank3[3913], bank2[3913], bank1[3913], bank0[3913]} = 32'h0;
    {bank3[3914], bank2[3914], bank1[3914], bank0[3914]} = 32'h0;
    {bank3[3915], bank2[3915], bank1[3915], bank0[3915]} = 32'h0;
    {bank3[3916], bank2[3916], bank1[3916], bank0[3916]} = 32'h0;
    {bank3[3917], bank2[3917], bank1[3917], bank0[3917]} = 32'h0;
    {bank3[3918], bank2[3918], bank1[3918], bank0[3918]} = 32'h0;
    {bank3[3919], bank2[3919], bank1[3919], bank0[3919]} = 32'h0;
    {bank3[3920], bank2[3920], bank1[3920], bank0[3920]} = 32'h0;
    {bank3[3921], bank2[3921], bank1[3921], bank0[3921]} = 32'h0;
    {bank3[3922], bank2[3922], bank1[3922], bank0[3922]} = 32'h0;
    {bank3[3923], bank2[3923], bank1[3923], bank0[3923]} = 32'h0;
    {bank3[3924], bank2[3924], bank1[3924], bank0[3924]} = 32'h0;
    {bank3[3925], bank2[3925], bank1[3925], bank0[3925]} = 32'h0;
    {bank3[3926], bank2[3926], bank1[3926], bank0[3926]} = 32'h0;
    {bank3[3927], bank2[3927], bank1[3927], bank0[3927]} = 32'h0;
    {bank3[3928], bank2[3928], bank1[3928], bank0[3928]} = 32'h0;
    {bank3[3929], bank2[3929], bank1[3929], bank0[3929]} = 32'h0;
    {bank3[3930], bank2[3930], bank1[3930], bank0[3930]} = 32'h0;
    {bank3[3931], bank2[3931], bank1[3931], bank0[3931]} = 32'h0;
    {bank3[3932], bank2[3932], bank1[3932], bank0[3932]} = 32'h0;
    {bank3[3933], bank2[3933], bank1[3933], bank0[3933]} = 32'h0;
    {bank3[3934], bank2[3934], bank1[3934], bank0[3934]} = 32'h0;
    {bank3[3935], bank2[3935], bank1[3935], bank0[3935]} = 32'h0;
    {bank3[3936], bank2[3936], bank1[3936], bank0[3936]} = 32'h0;
    {bank3[3937], bank2[3937], bank1[3937], bank0[3937]} = 32'h0;
    {bank3[3938], bank2[3938], bank1[3938], bank0[3938]} = 32'h0;
    {bank3[3939], bank2[3939], bank1[3939], bank0[3939]} = 32'h0;
    {bank3[3940], bank2[3940], bank1[3940], bank0[3940]} = 32'h0;
    {bank3[3941], bank2[3941], bank1[3941], bank0[3941]} = 32'h0;
    {bank3[3942], bank2[3942], bank1[3942], bank0[3942]} = 32'h0;
    {bank3[3943], bank2[3943], bank1[3943], bank0[3943]} = 32'h0;
    {bank3[3944], bank2[3944], bank1[3944], bank0[3944]} = 32'h0;
    {bank3[3945], bank2[3945], bank1[3945], bank0[3945]} = 32'h0;
    {bank3[3946], bank2[3946], bank1[3946], bank0[3946]} = 32'h0;
    {bank3[3947], bank2[3947], bank1[3947], bank0[3947]} = 32'h0;
    {bank3[3948], bank2[3948], bank1[3948], bank0[3948]} = 32'h0;
    {bank3[3949], bank2[3949], bank1[3949], bank0[3949]} = 32'h0;
    {bank3[3950], bank2[3950], bank1[3950], bank0[3950]} = 32'h0;
    {bank3[3951], bank2[3951], bank1[3951], bank0[3951]} = 32'h0;
    {bank3[3952], bank2[3952], bank1[3952], bank0[3952]} = 32'h0;
    {bank3[3953], bank2[3953], bank1[3953], bank0[3953]} = 32'h0;
    {bank3[3954], bank2[3954], bank1[3954], bank0[3954]} = 32'h0;
    {bank3[3955], bank2[3955], bank1[3955], bank0[3955]} = 32'h0;
    {bank3[3956], bank2[3956], bank1[3956], bank0[3956]} = 32'h0;
    {bank3[3957], bank2[3957], bank1[3957], bank0[3957]} = 32'h0;
    {bank3[3958], bank2[3958], bank1[3958], bank0[3958]} = 32'h0;
    {bank3[3959], bank2[3959], bank1[3959], bank0[3959]} = 32'h0;
    {bank3[3960], bank2[3960], bank1[3960], bank0[3960]} = 32'h0;
    {bank3[3961], bank2[3961], bank1[3961], bank0[3961]} = 32'h0;
    {bank3[3962], bank2[3962], bank1[3962], bank0[3962]} = 32'h0;
    {bank3[3963], bank2[3963], bank1[3963], bank0[3963]} = 32'h0;
    {bank3[3964], bank2[3964], bank1[3964], bank0[3964]} = 32'h0;
    {bank3[3965], bank2[3965], bank1[3965], bank0[3965]} = 32'h0;
    {bank3[3966], bank2[3966], bank1[3966], bank0[3966]} = 32'h0;
    {bank3[3967], bank2[3967], bank1[3967], bank0[3967]} = 32'h0;
    {bank3[3968], bank2[3968], bank1[3968], bank0[3968]} = 32'h0;
    {bank3[3969], bank2[3969], bank1[3969], bank0[3969]} = 32'h0;
    {bank3[3970], bank2[3970], bank1[3970], bank0[3970]} = 32'h0;
    {bank3[3971], bank2[3971], bank1[3971], bank0[3971]} = 32'h0;
    {bank3[3972], bank2[3972], bank1[3972], bank0[3972]} = 32'h0;
    {bank3[3973], bank2[3973], bank1[3973], bank0[3973]} = 32'h0;
    {bank3[3974], bank2[3974], bank1[3974], bank0[3974]} = 32'h0;
    {bank3[3975], bank2[3975], bank1[3975], bank0[3975]} = 32'h0;
    {bank3[3976], bank2[3976], bank1[3976], bank0[3976]} = 32'h0;
    {bank3[3977], bank2[3977], bank1[3977], bank0[3977]} = 32'h0;
    {bank3[3978], bank2[3978], bank1[3978], bank0[3978]} = 32'h0;
    {bank3[3979], bank2[3979], bank1[3979], bank0[3979]} = 32'h0;
    {bank3[3980], bank2[3980], bank1[3980], bank0[3980]} = 32'h0;
    {bank3[3981], bank2[3981], bank1[3981], bank0[3981]} = 32'h0;
    {bank3[3982], bank2[3982], bank1[3982], bank0[3982]} = 32'h0;
    {bank3[3983], bank2[3983], bank1[3983], bank0[3983]} = 32'h0;
    {bank3[3984], bank2[3984], bank1[3984], bank0[3984]} = 32'h0;
    {bank3[3985], bank2[3985], bank1[3985], bank0[3985]} = 32'h0;
    {bank3[3986], bank2[3986], bank1[3986], bank0[3986]} = 32'h0;
    {bank3[3987], bank2[3987], bank1[3987], bank0[3987]} = 32'h0;
    {bank3[3988], bank2[3988], bank1[3988], bank0[3988]} = 32'h0;
    {bank3[3989], bank2[3989], bank1[3989], bank0[3989]} = 32'h0;
    {bank3[3990], bank2[3990], bank1[3990], bank0[3990]} = 32'h0;
    {bank3[3991], bank2[3991], bank1[3991], bank0[3991]} = 32'h0;
    {bank3[3992], bank2[3992], bank1[3992], bank0[3992]} = 32'h0;
    {bank3[3993], bank2[3993], bank1[3993], bank0[3993]} = 32'h0;
    {bank3[3994], bank2[3994], bank1[3994], bank0[3994]} = 32'h0;
    {bank3[3995], bank2[3995], bank1[3995], bank0[3995]} = 32'h0;
    {bank3[3996], bank2[3996], bank1[3996], bank0[3996]} = 32'h0;
    {bank3[3997], bank2[3997], bank1[3997], bank0[3997]} = 32'h0;
    {bank3[3998], bank2[3998], bank1[3998], bank0[3998]} = 32'h0;
    {bank3[3999], bank2[3999], bank1[3999], bank0[3999]} = 32'h0;
    {bank3[4000], bank2[4000], bank1[4000], bank0[4000]} = 32'h0;
    {bank3[4001], bank2[4001], bank1[4001], bank0[4001]} = 32'h0;
    {bank3[4002], bank2[4002], bank1[4002], bank0[4002]} = 32'h0;
    {bank3[4003], bank2[4003], bank1[4003], bank0[4003]} = 32'h0;
    {bank3[4004], bank2[4004], bank1[4004], bank0[4004]} = 32'h0;
    {bank3[4005], bank2[4005], bank1[4005], bank0[4005]} = 32'h0;
    {bank3[4006], bank2[4006], bank1[4006], bank0[4006]} = 32'h0;
    {bank3[4007], bank2[4007], bank1[4007], bank0[4007]} = 32'h0;
    {bank3[4008], bank2[4008], bank1[4008], bank0[4008]} = 32'h0;
    {bank3[4009], bank2[4009], bank1[4009], bank0[4009]} = 32'h0;
    {bank3[4010], bank2[4010], bank1[4010], bank0[4010]} = 32'h0;
    {bank3[4011], bank2[4011], bank1[4011], bank0[4011]} = 32'h0;
    {bank3[4012], bank2[4012], bank1[4012], bank0[4012]} = 32'h0;
    {bank3[4013], bank2[4013], bank1[4013], bank0[4013]} = 32'h0;
    {bank3[4014], bank2[4014], bank1[4014], bank0[4014]} = 32'h0;
    {bank3[4015], bank2[4015], bank1[4015], bank0[4015]} = 32'h0;
    {bank3[4016], bank2[4016], bank1[4016], bank0[4016]} = 32'h0;
    {bank3[4017], bank2[4017], bank1[4017], bank0[4017]} = 32'h0;
    {bank3[4018], bank2[4018], bank1[4018], bank0[4018]} = 32'h0;
    {bank3[4019], bank2[4019], bank1[4019], bank0[4019]} = 32'h0;
    {bank3[4020], bank2[4020], bank1[4020], bank0[4020]} = 32'h0;
    {bank3[4021], bank2[4021], bank1[4021], bank0[4021]} = 32'h0;
    {bank3[4022], bank2[4022], bank1[4022], bank0[4022]} = 32'h0;
    {bank3[4023], bank2[4023], bank1[4023], bank0[4023]} = 32'h0;
    {bank3[4024], bank2[4024], bank1[4024], bank0[4024]} = 32'h0;
    {bank3[4025], bank2[4025], bank1[4025], bank0[4025]} = 32'h0;
    {bank3[4026], bank2[4026], bank1[4026], bank0[4026]} = 32'h0;
    {bank3[4027], bank2[4027], bank1[4027], bank0[4027]} = 32'h0;
    {bank3[4028], bank2[4028], bank1[4028], bank0[4028]} = 32'h0;
    {bank3[4029], bank2[4029], bank1[4029], bank0[4029]} = 32'h0;
    {bank3[4030], bank2[4030], bank1[4030], bank0[4030]} = 32'h0;
    {bank3[4031], bank2[4031], bank1[4031], bank0[4031]} = 32'h0;
    {bank3[4032], bank2[4032], bank1[4032], bank0[4032]} = 32'h0;
    {bank3[4033], bank2[4033], bank1[4033], bank0[4033]} = 32'h0;
    {bank3[4034], bank2[4034], bank1[4034], bank0[4034]} = 32'h0;
    {bank3[4035], bank2[4035], bank1[4035], bank0[4035]} = 32'h0;
    {bank3[4036], bank2[4036], bank1[4036], bank0[4036]} = 32'h0;
    {bank3[4037], bank2[4037], bank1[4037], bank0[4037]} = 32'h0;
    {bank3[4038], bank2[4038], bank1[4038], bank0[4038]} = 32'h0;
    {bank3[4039], bank2[4039], bank1[4039], bank0[4039]} = 32'h0;
    {bank3[4040], bank2[4040], bank1[4040], bank0[4040]} = 32'h0;
    {bank3[4041], bank2[4041], bank1[4041], bank0[4041]} = 32'h0;
    {bank3[4042], bank2[4042], bank1[4042], bank0[4042]} = 32'h0;
    {bank3[4043], bank2[4043], bank1[4043], bank0[4043]} = 32'h0;
    {bank3[4044], bank2[4044], bank1[4044], bank0[4044]} = 32'h0;
    {bank3[4045], bank2[4045], bank1[4045], bank0[4045]} = 32'h0;
    {bank3[4046], bank2[4046], bank1[4046], bank0[4046]} = 32'h0;
    {bank3[4047], bank2[4047], bank1[4047], bank0[4047]} = 32'h0;
    {bank3[4048], bank2[4048], bank1[4048], bank0[4048]} = 32'h0;
    {bank3[4049], bank2[4049], bank1[4049], bank0[4049]} = 32'h0;
    {bank3[4050], bank2[4050], bank1[4050], bank0[4050]} = 32'h0;
    {bank3[4051], bank2[4051], bank1[4051], bank0[4051]} = 32'h0;
    {bank3[4052], bank2[4052], bank1[4052], bank0[4052]} = 32'h0;
    {bank3[4053], bank2[4053], bank1[4053], bank0[4053]} = 32'h0;
    {bank3[4054], bank2[4054], bank1[4054], bank0[4054]} = 32'h0;
    {bank3[4055], bank2[4055], bank1[4055], bank0[4055]} = 32'h0;
    {bank3[4056], bank2[4056], bank1[4056], bank0[4056]} = 32'h0;
    {bank3[4057], bank2[4057], bank1[4057], bank0[4057]} = 32'h0;
    {bank3[4058], bank2[4058], bank1[4058], bank0[4058]} = 32'h0;
    {bank3[4059], bank2[4059], bank1[4059], bank0[4059]} = 32'h0;
    {bank3[4060], bank2[4060], bank1[4060], bank0[4060]} = 32'h0;
    {bank3[4061], bank2[4061], bank1[4061], bank0[4061]} = 32'h0;
    {bank3[4062], bank2[4062], bank1[4062], bank0[4062]} = 32'h0;
    {bank3[4063], bank2[4063], bank1[4063], bank0[4063]} = 32'h0;
    {bank3[4064], bank2[4064], bank1[4064], bank0[4064]} = 32'h0;
    {bank3[4065], bank2[4065], bank1[4065], bank0[4065]} = 32'h0;
    {bank3[4066], bank2[4066], bank1[4066], bank0[4066]} = 32'h0;
    {bank3[4067], bank2[4067], bank1[4067], bank0[4067]} = 32'h0;
    {bank3[4068], bank2[4068], bank1[4068], bank0[4068]} = 32'h0;
    {bank3[4069], bank2[4069], bank1[4069], bank0[4069]} = 32'h0;
    {bank3[4070], bank2[4070], bank1[4070], bank0[4070]} = 32'h0;
    {bank3[4071], bank2[4071], bank1[4071], bank0[4071]} = 32'h0;
    {bank3[4072], bank2[4072], bank1[4072], bank0[4072]} = 32'h0;
    {bank3[4073], bank2[4073], bank1[4073], bank0[4073]} = 32'h0;
    {bank3[4074], bank2[4074], bank1[4074], bank0[4074]} = 32'h0;
    {bank3[4075], bank2[4075], bank1[4075], bank0[4075]} = 32'h0;
    {bank3[4076], bank2[4076], bank1[4076], bank0[4076]} = 32'h0;
    {bank3[4077], bank2[4077], bank1[4077], bank0[4077]} = 32'h0;
    {bank3[4078], bank2[4078], bank1[4078], bank0[4078]} = 32'h0;
    {bank3[4079], bank2[4079], bank1[4079], bank0[4079]} = 32'h0;
    {bank3[4080], bank2[4080], bank1[4080], bank0[4080]} = 32'h0;
    {bank3[4081], bank2[4081], bank1[4081], bank0[4081]} = 32'h0;
    {bank3[4082], bank2[4082], bank1[4082], bank0[4082]} = 32'h0;
    {bank3[4083], bank2[4083], bank1[4083], bank0[4083]} = 32'h0;
    {bank3[4084], bank2[4084], bank1[4084], bank0[4084]} = 32'h0;
    {bank3[4085], bank2[4085], bank1[4085], bank0[4085]} = 32'h0;
    {bank3[4086], bank2[4086], bank1[4086], bank0[4086]} = 32'h0;
    {bank3[4087], bank2[4087], bank1[4087], bank0[4087]} = 32'h0;
    {bank3[4088], bank2[4088], bank1[4088], bank0[4088]} = 32'h0;
    {bank3[4089], bank2[4089], bank1[4089], bank0[4089]} = 32'h0;
    {bank3[4090], bank2[4090], bank1[4090], bank0[4090]} = 32'h0;
    {bank3[4091], bank2[4091], bank1[4091], bank0[4091]} = 32'h0;
    {bank3[4092], bank2[4092], bank1[4092], bank0[4092]} = 32'h0;
    {bank3[4093], bank2[4093], bank1[4093], bank0[4093]} = 32'h0;
    {bank3[4094], bank2[4094], bank1[4094], bank0[4094]} = 32'h0;
    {bank3[4095], bank2[4095], bank1[4095], bank0[4095]} = 32'h0;


     end

endmodule
